.option geoshrink=0.9
.param ccoflag=0 rgflag=0 sigma_factor=1 rcoflag=0 scale_mos=0.9 designflag_mos=0 bidirectionflag_mos=1 iboffn_flag=0 totalflag_mos=1 globalflag_mos=1 mismatchflag_mos=1 global_factor=1 local_factor=1 iboffp_flag=0 noiseflagn=0 noiseflagp=0 noiseflagn_mc=0 noiseflagp_mc=0 sigma_factor_flicker=1
.param toxn=1.95e-009                dxln=0                        dxwn=0 cjn=1.428e-03                cjswn=1.069e-10                cjswgn=2.9e-10 cgon=8.14e-011                cgln=2.4209e-011              ddlcn='5.81e-009-(5.81e-009)' cfn='6.62e-011+9.73e-11*ccoflag' ntoxn=1 dvthn=0                        dlvthn=0                        dwvthn=0 dpvthn=0                        du0n=0                        dlu0n=0 dwu0n=0                        dpu0n=0                        dvsatn=0 dlvsatn=0                        dwvsatn=0                        dpvsatn=0 dk2n=0                        dlk2n=0                        dwk2n=0 dpk2n=0                        dvoffn=0                        dlvoffn=0 dwvoffn=0                        dpvoffn=0                        dpdiblc2n=0 dlpdiblc2n=0                        dwpdiblc2n=0                        dppdiblc2n=0 dagsn=0                        dlagsn=0                        dwagsn=0 dpagsn=0                        dnfactorn=0                        dlnfactorn=0 dwnfactorn=0                        dpnfactorn=0                        dcitn=0 dlcitn=0                        dwcitn=0                        dpcitn=0 deta0n=0                        dleta0n=0                        dweta0n=0 dpeta0n=0                        dpclmn=0                        dlpclmn=0 dwpclmn=0                        dppclmn=0                        jtsswgn='4.52e-005*(1+1.57*iboffn_flag)' dminvn=0                        dketan=0                        dlketan=0 dwketan=0                        dpketan=0                        dua1n=0 dlua1n=0                        dwua1n=0                        dpua1n=0 datn=0                        dlatn=0                        dwatn=0 dpatn=0 ss_flagn=0                        ff_flagn=0                        sf_flagn=0                        fs_flagn=0 monte_flagn=0
.param toxp=2.18e-009                dxlp=0                        dxwp=0 cjp=1.514e-03                cjswp=1.129e-10                cjswgp=2.08e-10 cgop=5.02e-011                cglp=6.0796e-011              ddlcp='6.67e-009-(6.67e-009)' cfp='9e-011+0.92e-10*ccoflag' ntoxp=1 dvthp=0                        dlvthp=0                        dwvthp=0 dpvthp=0                        dk2p=0                        dlk2p=0 dwk2p=0                        dpk2p=0                        deta0p=0 dleta0p=0                        dweta0p=0                        dpeta0p=0 dvoffp=0                        dlvoffp=0                        dwvoffp=0 dpvoffp=0                        dcitp=0                        dlcitp=0 dwcitp=0                        dpcitp=0                        dnfactorp=0 dlnfactorp=0                        dwnfactorp=0                        dpnfactorp=0 du0p=0                        dlu0p=0                        dwu0p=0 dpu0p=0                        dpclmp=0                        dlpclmp=0 dwpclmp=0                        dppclmp=0                        dpdiblc2p=0 dlpdiblc2p=0                        dvsatp=0                        dlvsatp=0 dwvsatp=0                        dpvsatp=0                        da0p=0 dagsp=0                        dwagsp=0                        dlagsp=0 dpagsp=0                        jtsswgp='1.5e-007*(1+0.55*iboffp_flag)' dminvp=0 datp=0                        dlatp=0                        dwatp=0 dpatp=0                        dua1p=0                        dlua1p=0 dwua1p=0                        dpua1p=0                        dketap=0 dlketap=0                        dwketap=0                        dpketap=0 ss_flagp=0                        ff_flagp=0                        sf_flagp=0                        fs_flagp=0 monte_flagp=0 c1fn=6.310000e+41             c2fn=1.380000e+24             c3fn=4.540000e+05 c1fp=2.200000e+41             c2fp=3.000000e+27             c3fp=1.000000e+11
.param ccoflag_12=0 rgflag_12=0 sigma_factor_12=1 rcoflag_12=0 scale_mos_12=0.9 iboffn_flag_12=0 iboffp_flag_12=0 totalflag_mos_12=1 globalflag_mos_12=1 mismatchflag_mos_12=1 global_factor_12=0.96 local_factor_12=1 noiseflagn_12=0 noiseflagp_12=0 noiseflagn_12_mc=0 noiseflagp_12_mc=0 sigma_factor_flicker_12=1
.param toxn_12=2.42e-009                dxln_12=0                        dxwn_12=0 cjn_12=0.00144                  cjswn_12=1.1300e-10               cjswgn_12=2.7000e-10 cgon_12=1.0000e-10               cgln_12=5.0000e-12               ddlcn_12='7.50e-09-(7.50e-09)' ntoxn_12=1                        cfn_12='6.7e-011+9.3e-011*ccoflag_12' dvthn_12=0                        dlvthn_12=0                        dwvthn_12=0 dpvthn_12=0                        du0n_12=0                        dlu0n_12=0 dwu0n_12=0                        dpu0n_12=0                        dvsatn_12=0 dlvsatn_12=0                        dwvsatn_12=0                        dpvsatn_12=0 dk2n_12=0                        dlk2n_12=0                        dwk2n_12=0 dpk2n_12=0                        dagsn_12=0                        dlagsn_12=0 dwagsn_12=0                        dpagsn_12=0                        dcitn_12=0 dlcitn_12=0                        dwcitn_12=0                        dpcitn_12=0 dpclmn_12=0                        dlpclmn_12=0                        dwpclmn_12=0 dppclmn_12=0                        dua1n_12=0                        dlua1n_12=0 dwua1n_12=0                        dpua1n_12=0                        ducn_12=0 dlucn_12=0                        dwucn_12=0                        dpucn_12=0 dketan_12=0                        dlketan_12=0                        dwketan_12=0 dpketan_12=0                        jtsswgn_12='2e-007*(1+21*0.3*iboffn_flag_12)' ss_flagn_12=0 ff_flagn_12=0 sf_flagn_12=0 fs_flagn_12=0 monte_flagn_12=0
.param toxp_12=2.687e-009               dxlp_12=0                        dxwp_12=0 cjp_12=0.001878                 cjswp_12=1.13e-10                 cjswgp_12=1.86e-10 cgop_12=9.20e-11                 cglp_12=1.00e-11                 ddlcp_12='8.00e-09-(8.00e-09)' ntoxp_12=1                        cfp_12='9.1e-011+8.7e-11*ccoflag_12' dvthp_12=0                        dlvthp_12=0                        dwvthp_12=0 dpvthp_12=0                        du0p_12=0                        dlu0p_12=0 dwu0p_12=0                        dpu0p_12=0                        dvsatp_12=0 dlvsatp_12=0                        dwvsatp_12=0                        dpvsatp_12=0 dk2p_12=0                        dlk2p_12=0                        dwk2p_12=0 dpk2p_12=0                        dvoffp_12=0                        dlvoffp_12=0 dwvoffp_12=0                        dpvoffp_12=0                        dagsp_12=0 dlagsp_12=0                        dwagsp_12=0                        dpagsp_12=0 dcitp_12=0                        dlcitp_12=0                        dwcitp_12=0 dpcitp_12=0                        deta0p_12=0                        dpclmp_12=0 dua1p_12=0                        dlua1p_12=0                        dwua1p_12=0 dpua1p_12=0                        ducp_12=0                        dlucp_12=0 dwucp_12=0                        dpucp_12=0                        dketap_12=0 dlketap_12=0                        dwketap_12=0                        dpketap_12=0 jtsswgp_12='1e-009*(1+1200*0.06*iboffp_flag_12)' ss_flagp_12=0 ff_flagp_12=0 sf_flagp_12=0 fs_flagp_12=0 monte_flagp_12=0 c1fn_12=7e+041                   c2fn_12=1e+023                   c3fn_12=1e+007 c1fp_12=1e+042                   c2fp_12=1e+027                   c3fp_12=6e+009
.param ccoflag_18=0 rgflag_18=0 sigma_factor_18=1 rcoflag_18=0 scale_mos_18=0.9 totalflag_mos_18=1 globalflag_mos_18=1 mismatchflag_mos_18=1 global_factor_18=1 local_factor_18=1 noiseflagn_18=0 noiseflagp_18=0 noiseflagn_18_mc=0 noiseflagp_18_mc=0 sigma_factor_flicker_18=1
.param toxn_18=3.36e-009                dxln_18=0                        dxwn_18=0 ddlcn_18='1.17e-008-(1.17e-008)'  cgon_18=4.50e-11                 cgln_18=7.90e-11 cjn_18=0.001472                 cjswn_18=1.086e-10                cjswgn_18=2.016e-10 cfn_18='8.09e-011+5.742e-11*ccoflag_18' dvthn_18=0 dwvthn_18=0                        dlvthn_18=0                        dpvthn_18=0 du0n_18=0                        dwu0n_18=0                        dlu0n_18=0 dpu0n_18=0                        dk2n_18=0                        dwk2n_18=0 dlk2n_18=0                        dpk2n_18=0                        dagsn_18=0 dwagsn_18=0                        dpdiblc2n_18=0                        dlpdiblc2n_18=0 dvsatn_18=0                        dwvsatn_18=0                        ducn_18=0 dlucn_18=0                        dwucn_18=0                        dpucn_18=0 dketan_18=0                        dlketan_18=0                        dwketan_18=0 dpketan_18=0
.param toxp_18=3.65e-009                dxlp_18=0                        dxwp_18=0 ddlcp_18='1.24e-008-(1.24e-008)'  cgop_18=7.5e-12                  cglp_18=1.105e-10 cjp_18=0.001836                 cjswp_18=1.454e-010               cjswgp_18=1.847e-10 cfp_18='9.43e-011+5.68e-11*ccoflag_18' dvthp_18=0 dwvthp_18=0                        dlvthp_18=0                        dpvthp_18=0 du0p_18=0                        dwu0p_18=0                        dlu0p_18=0 dpu0p_18=0                        dk2p_18=0                        dwk2p_18=0 dlk2p_18=0                        dpk2p_18=0                        dagsp_18=0 dwagsp_18=0                        dpdiblc2p_18=0                        dlpdiblc2p_18=0 dvsatp_18=0                        dwvsatp_18=0                        ducp_18=0 dlucp_18=0                        dwucp_18=0                        dpucp_18=0 dvoffp_18=0                        dlvoffp_18=0                        dwvoffp_18=0 dpvoffp_18=0                        dpkt1p_18=0                        dltvoffp_18=0 dkt2p_18=0                        duc1p_18=0                        dlub1p_18=0 dlketap_18=0 ss_flagp_18=0 ff_flagp_18=0 sf_flagp_18=0 fs_flagp_18=0 monte_flagn_18=0 monte_flagp_18=0 c1fn_18=2.31e+041                c2fn_18=1.18e+022                c3fn_18=1.44e+008 c1fp_18=3.56e+041                c2fp_18=4.89e+026                c3fp_18=5.92e+005
.param ccoflag_18ud15=0 rgflag_18ud15=0 sigma_factor_18ud15=1 rcoflag_18ud15=0 scale_mos_18ud15=0.9 totalflag_mos_18ud15=1 globalflag_mos_18ud15=1 mismatchflag_mos_18ud15=1 global_factor_18ud15=1 local_factor_18ud15=1 noiseflagn_18ud15=0 noiseflagp_18ud15=0 noiseflagn_18ud15_mc=0 noiseflagp_18ud15_mc=0 sigma_factor_flicker_18ud15=1
.param toxn_18ud15=3.36e-009                dxln_18ud15=0                        dxwn_18ud15=0 ddlcn_18ud15='1.17e-008-(1.17e-008)'  cgon_18ud15=4.50e-11                 cgln_18ud15=7.90e-11 cjn_18ud15=0.001472                 cjswn_18ud15=1.086e-10                cjswgn_18ud15=2.016e-10 cfn_18ud15='8.09e-011+5.742e-11*ccoflag_18ud15' dvthn_18ud15=0 dwvthn_18ud15=0                        dlvthn_18ud15=0                        dpvthn_18ud15=0 du0n_18ud15=0                        dwu0n_18ud15=0                        dlu0n_18ud15=0 dpu0n_18ud15=0                        dk2n_18ud15=0                        dwk2n_18ud15=0 dlk2n_18ud15=0                        dpk2n_18ud15=0                        dagsn_18ud15=0 dwagsn_18ud15=0                        dpdiblc2n_18ud15=0                        dlpdiblc2n_18ud15=0 dvsatn_18ud15=0                        dwvsatn_18ud15=0                        ducn_18ud15=0 dlucn_18ud15=0                        dwucn_18ud15=0                        dpucn_18ud15=0 dketan_18ud15=0                        dlketan_18ud15=0                        dwketan_18ud15=0 dpketan_18ud15=0
.param toxp_18ud15=3.65e-009                dxlp_18ud15=0                        dxwp_18ud15=0 ddlcp_18ud15='1.24e-008-(1.24e-008)'  cgop_18ud15=7.5e-12                  cglp_18ud15=1.105e-10 cjp_18ud15=0.001836                 cjswp_18ud15=1.454e-010               cjswgp_18ud15=1.847e-10 cfp_18ud15='9.43e-011+5.68e-11*ccoflag_18ud15' dvthp_18ud15=0 dwvthp_18ud15=0                        dlvthp_18ud15=0                        dpvthp_18ud15=0 du0p_18ud15=0                        dwu0p_18ud15=0                        dlu0p_18ud15=0 dpu0p_18ud15=0                        dk2p_18ud15=0                        dwk2p_18ud15=0 dlk2p_18ud15=0                        dpk2p_18ud15=0                        dagsp_18ud15=0 dwagsp_18ud15=0                        dpdiblc2p_18ud15=0                        dlpdiblc2p_18ud15=0 dvsatp_18ud15=0                        dwvsatp_18ud15=0                        ducp_18ud15=0 dlucp_18ud15=0                        dwucp_18ud15=0                        dpucp_18ud15=0 dvoffp_18ud15=0                        dlvoffp_18ud15=0                        dwvoffp_18ud15=0 dpvoffp_18ud15=0                        dpkt1p_18ud15=0                        dltvoffp_18ud15=0 dkt2p_18ud15=0                        duc1p_18ud15=0                        dlub1p_18ud15=0 dlketap_18ud15=0 ss_flagp_18ud15=0 ff_flagp_18ud15=0 sf_flagp_18ud15=0 fs_flagp_18ud15=0 monte_flagn_18ud15=0 monte_flagp_18ud15=0 c1fn_18ud15=2.31e+041                c2fn_18ud15=1.18e+022                c3fn_18ud15=1.44e+008 c1fp_18ud15=3.56e+041                c2fp_18ud15=4.89e+026                c3fp_18ud15=5.92e+005
.param ccoflag_hia=0 rgflag_hia=0 sigma_factor_hia=1 iboffn_flag_hia=0 rcoflag_hia=0 scale_mos_hia=0.9
.param toxn_hia=1.95e-009                dxln_hia=0                        dxwn_hia=0 cjn_hia=1.428e-03                cjswn_hia=1.069e-10                cjswgn_hia=2.9e-10 cgon_hia=8.14e-011                cgln_hia=2.4209e-011              ddlcn_hia='5.81e-009-(5.81e-009)' cfn_hia='6.62e-011+9.73e-11*ccoflag_hia' ntoxn_hia=1 dvthn_hia=0                        dlvthn_hia=0                        dwvthn_hia=0 dpvthn_hia=0                        du0n_hia=0                        dlu0n_hia=0 dwu0n_hia=0                        dpu0n_hia=0                        dubn_hia=0 dlubn_hia=0                        dwubn_hia=0                        dpubn_hia=0 dvsatn_hia=0                        dlvsatn_hia=0                        dwvsatn_hia=0 dpvsatn_hia=0                        dk2n_hia=0                        dlk2n_hia=0 dwk2n_hia=0                        dpk2n_hia=0                        dvoffn_hia=0 dlvoffn_hia=0                        dwvoffn_hia=0                        dpvoffn_hia=0 dpdiblc2n_hia=0                        dlpdiblc2n_hia=0                        dwpdiblc2n_hia=0 dppdiblc2n_hia=0                        da0n_hia=0                        dla0n_hia=0 dwa0n_hia=0                        dpa0n_hia=0                        dagsn_hia=0 dlagsn_hia=0                        dwagsn_hia=0                        dpagsn_hia=0 dnfactorn_hia=0                        dlnfactorn_hia=0                        dwnfactorn_hia=0 dpnfactorn_hia=0                        dcitn_hia=0                        dlcitn_hia=0 dwcitn_hia=0                        dpcitn_hia=0                        deta0n_hia=0 dleta0n_hia=0                        dweta0n_hia=0                        dpeta0n_hia=0 dpclmn_hia=0                        dlpclmn_hia=0                        dwpclmn_hia=0 dppclmn_hia=0                        jtsswgn_hia='4.52e-005*(1+1.57*iboffn_flag_hia)' dminvn_hia=0 dketan_hia=0                        dlketan_hia=0                        dwketan_hia=0 dpketan_hia=0                        dua1n_hia=0                        dlua1n_hia=0 dwua1n_hia=0                        dpua1n_hia=0                        datn_hia=0 dlatn_hia=0                        dwatn_hia=0                        dpatn_hia=0
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_hia_mac.global nmos ( modelid=17                         level=54                         lmin=0.09e-06 lmax=0.13601e-6                 wmin=13.5e-06                   wmax=54.01e-06 version=4.5                        binunit=2                          paramchk=1 mobmod=0                          capmod=2                          igcmod=1 igbmod=1                          diomod=1                          rdsmod=0 rbodymod=0                          rgatemod='1*rgflag_hia'             permod=1 acnqsmod=0                          trnqsmod=0                          tempmod=0 tnom=25                         toxe=1.95e-009                  toxm=1.95e-009 dtox=4.06e-010                  epsrox=3.9                        wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=-4e-009 xw=6e-009                     dlc=5.81e-009                  dwc=0 xpart=1                          toxref=3e-009                     dlcig=2.5e-009 vth0=0.36964921                 lvth0=-2.1198317e-009            k1=0.3372 k2=-0.013473796               lk2=1.5499559e-010             k3=-1 k3b=0.8                        w0=0                          dvt0=0.88 dvt1=0.79                       dvt2=0.48                       dvt0w=0 dvt1w=0                          dvt2w=0                          dsub=0.6 minv=-0.42453                   voffl=0                          dvtp0=1e-006 dvtp1=1.4                        lpe0=0                          lpeb=0 xj=6.7e-008                   ngate=1.476e+020                 ndep=1e+017 nsd=1e+020                     phin=0.13375                    cdsc=0 cdscb=0                          cdscd=0                          cit=0.0014925714 lcit=2.1357486e-010             voff=-0.18155479                lvoff=-1.9302884e-009 nfactor=0.7                        eta0=0.009                      etab=-0.035607824 letab=-1.4469841e-016            ud=0                          lud=0 wud=0                          pud=0                          u0=0.023679413 lu0=-4.6563949e-010            ua=-1.555546e-009             lua=-1.3558241e-017 ub=2.0010159e-018             lub=-2.1415365e-026            uc=1.2501587e-010 luc=-3.1833651e-018            vsat=88841.27                   lvsat=0.0044856508 a0=2.9555556                  la0=-2.0257778e-007            ags=4.952381 lags=4.3409524e-007             a1=0                          a2=1 b0=0                          b1=0                          keta=-0.061746032 lketa=-1.4469841e-008            dwg=0                          dwb=0 pclm=0.93171238                 lpclm=1.4472735e-008             pdiblc1=0 pdiblc2=0.003                      pdiblcb=1                          drout=0.56 pvag=2                          delta=0.01                       pscbe1=1e+009 pscbe2=1e-020                     fprout=78                         pdits=0.0027 pditsd=0                          pditsl=0                          rsh=18.0 rdsw=120                        rsw=0                          rdw=0 prwg=0                          prwb=0                          wr=1 alpha0=1e-008                     alpha1=1.5                        beta0=12 agidl=1e-006                     bgidl=3.459e+009                 cgidl=0.295 egidl=0.27814                    aigbacc=0.013638318                laigbacc=-9.1015302e-011 bigbacc=0.0074708                  cigbacc=0.2809                     nigbacc=4.05 aigbinv=0.2415                     bigbinv=0.0309                     cigbinv=0.006 eigbinv=1.1                        nigbinv=1                          aigc=0.010861235 laigc=-1.037806e-011             bigc=0.00159                    cigc=1e-005 aigsd=0.0097591825               laigsd=-9.2606984e-012            bigsd=0.00041057365 lbigsd=8.019186e-012              cigsd=2e-020                     nigc=3.083 poxedge=1                          pigcd=2.46                       ntox=1 xrcrg1=12                         xrcrg2=1                          vfbsdoff=0.01 lvfbsdoff=0                          wvfbsdoff=0                          pvfbsdoff=0 cgso=8.14e-011                  cgdo=8.14e-011                  cgbo=0 cgdl=2.4209e-011                cgsl=2.4209e-011                clc=0 cle=0.6                        cf='6.62e-011+9.73e-11*ccoflag_hia' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=6.5                        noff=2.5                        voffcv=-0.098559 tvoff=0.00218524                 ltvoff=-2.39635e-011              wtvoff=0 ptvoff=0                          tvfbsdoff=0.1                        ltvfbsdoff=0 wtvfbsdoff=0                          ptvfbsdoff=0                          kt1=-0.16675705 lkt1=-2.4119692e-009            kt1l=0                          kt2=-0.073319397 lkt2=1.9210161e-009             ute=-1                         ua1=1.2818459e-009 lua1=-9.9995285e-017            ub1=-1.3452089e-018            lub1=1.0196752e-025 uc1=5.0920635e-011             luc1=-2.3151746e-018            prt=0 at=88395.067                  lat=-0.0017420426              fnoimod=1 tnoimod=0                          em=1e+006                     ef=0.9 noia=6.31e+041                  noib=1.38e+024                  noic=454000 lintnoi=-2.79e-008                 jss=4.32e-07                   jsd=4.32e-07 jsws=1.17e-13                   jswd=1.17e-13                   jswgs=1.17e-13 jswgd=1.17e-13                   njs=1.03                       njd=1.03 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=8.219999                   bvd=8.219999 xjbvs=1                          xjbvd=1                          njtsswg=16 xtsswgs=0.16                       xtsswgd=0.16                       tnjtsswg=1 vtsswgs=1                          vtsswgd=1                          pbs=0.672 pbd=0.672                      cjs=0.001428                   cjd=0.001428 mjs=0.321                      mjd=0.321                      pbsws=0.480 pbswd=0.480                      cjsws=1.069e-010                 cjswd=1.069e-010 mjsws=0.016                      mjswd=0.016                      pbswgs=0.990 pbswgd=0.990                      cjswgs=2.9e-010                   cjswgd=2.9e-010 mjswgs=0.725                      mjswgd=0.725                      tpb=0.00114 tcj=0.00072                    tpbsw=0.00244                    tcjsw=0.00020 tpbswg=0.00171                    tcjswg=0.00124                    xtis=3 xtid=3                          dmcg=3.8e-008                   dmci=3.8e-008 dmdg=0                          dmcgt=0                          dwj=0 xgw=0                          xgl=2.64e-009                  rshg=16.42 gbmin=1e-012                     rbpb=50                         rbpd=50 rbps=50                         rbdb=50                         rbsb=50 ngcon=1                          leta0=0                          lnfactor=0 lpdiblc2=0                          pa0=0                          pags=0 pat=0                          pcit=0                          peta0=0 pk2=0                          pketa=0                          pnfactor=0 ppclm=0                          ppdiblc2=0                          pu0=0 pua1=0                          pub=0                          pvoff=0 pvsat=0                          pvth0=0                          wa0=0 wags=0                          wat=0                          wcit=0 weta0=0                          wk2=0                          wketa=0 wnfactor=0                          wpclm=0                          wpdiblc2=0 wu0=0                          wua1=0                          wub=0 wvoff=0                          wvsat=0                          wvth0=0 pk2we=0                          lk2we=0                          wk2we=0 k2we=0.0000                     pku0we=-1e-18                     wku0we=3e-11 lku0we=4.5e-11                    ku0we=-0.0016                    pkvth0we=1.3e-018 wkvth0we=-4.1e-011                  lkvth0we=-1.05e-011                 kvth0we=0.00053 wec=-9093.6                    web=2153.1                     scref=1e-6 wpemod=1 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.2                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.0 tmi_ver_mcratio=0.0                    tmi_ver_mcglobal=0.0                   tmi_ver_mclocal=0.0 tmi_ver_mcdelta=0.0                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.0 iboffn_flag='iboffn_flag_hia' sigma_factor='sigma_factor_hia' ccoflag='ccoflag_hia' rcoflag='rcoflag_hia' rgflag='rgflag_hia' delvto=0 mulu0=1 dlc_fmt=2 tox_c='toxn_hia'                 dxl_c='dxln_hia'                 dxw_c='dxwn_hia' cj_c='cjn_hia'                  cjsw_c='cjswn_hia'                cjswg_c='cjswgn_hia' cgo_c='cgon_hia'                 cgl_c='cgln_hia'                 ddlc_c='ddlcn_hia' cf_c='cfn_hia'                  ntox_c='ntoxn_hia'                dvth_c='dvthn_hia' dlvth_c='dlvthn_hia'               dwvth_c='dwvthn_hia'               dpvth_c='dpvthn_hia' du0_c='du0n_hia'                 dlu0_c='dlu0n_hia'                dwu0_c='dwu0n_hia' dpu0_c='dpu0n_hia'                dub_c='dubn_hia'                 dlub_c='dlubn_hia' dwub_c='dwubn_hia'                dpub_c='dpubn_hia'                dvsat_c='dvsatn_hia' dlvsat_c='dlvsatn_hia'              dwvsat_c='dwvsatn_hia'              dpvsat_c='dpvsatn_hia' dk2_c='dk2n_hia'                 dlk2_c='dlk2n_hia'                dwk2_c='dwk2n_hia' dpk2_c='dpk2n_hia'                dvoff_c='dvoffn_hia'               dlvoff_c='dlvoffn_hia' dwvoff_c='dwvoffn_hia'              dpvoff_c='dpvoffn_hia'              dpdiblc2_c='dpdiblc2n_hia' dlpdiblc2_c='dlpdiblc2n_hia'           dwpdiblc2_c='dwpdiblc2n_hia'           dppdiblc2_c='dppdiblc2n_hia' da0_c='da0n_hia'                 dla0_c='dla0n_hia'                dwa0_c='dwa0n_hia' dpa0_c='dpa0n_hia'                dags_c='dagsn_hia'                dlags_c='dlagsn_hia' dwags_c='dwagsn_hia'               dpags_c='dpagsn_hia'               dnfactor_c='dnfactorn_hia' dlnfactor_c='dlnfactorn_hia'           dwnfactor_c='dwnfactorn_hia'           dpnfactor_c='dpnfactorn_hia' dcit_c='dcitn_hia'                dlcit_c='dlcitn_hia'               dwcit_c='dwcitn_hia' dpcit_c='dpcitn_hia'               deta0_c='deta0n_hia'               dleta0_c='dleta0n_hia' dweta0_c='dweta0n_hia'              dpeta0_c='dpeta0n_hia'              dpclm_c='dpclmn_hia' dlpclm_c='dlpclmn_hia'              dwpclm_c='dwpclmn_hia'              dppclm_c='dppclmn_hia' jtsswg_c='jtsswgn_hia'              dminv_c='dminvn_hia'               dketa_c='dketan_hia' dlketa_c='dlketan_hia'              dwketa_c='dwketan_hia'              dpketa_c='dpketan_hia' dua1_c='dua1n_hia'                dlua1_c='dlua1n_hia'               dwua1_c='dwua1n_hia' dpua1_c='dpua1n_hia'               dat_c='datn_hia'                 dlat_c='dlatn_hia' dwat_c='dwatn_hia'                dpat_c='dpatn_hia' xw0=6e-09                      xl0=-4e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0 cf0=6.62e-011                  cco=9.73e-11 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.49                       l_rjtsswg=2.5e-5                     ll_rjtsswg=3 w_rjtsswg=0                          ww_rjtsswg=0                          p_rjtsswg=0 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6                sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=0                   lreflod=1e-6                llodref=3 lod_clamp=-1e90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=1 kvth00=0                   lkvth00=0                   wkvth00=0 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=0                   lku000=0                   wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0                   lkvth000=0                   wkvth000=0         		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=0                   wku01=0 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=0                   wkvth01=0 pkvth01=0                   llodvth1=1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.06               lku02=1.5e-7              wku02=7e-8 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=-0.5 kvth02=7e-3                lkvth02=-9e-9               wkvth02=16e-9 pkvth02=1e-15               llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=-0.03               lku03=7e5                 wku03=-5e-8 pku03=0                   tku03=0                   llodku03=-1 wlodku03=1                   kvsat3=0 kvth03=9e-3                lkvth03=-3e-9               wkvth03=-2e-8 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=-0.000                   lku003=-0.0e-9                   wku003=-0e-9         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0.0e-3                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='0.15*01'           wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl='1.4e-12*1'         ldplkvth0=1.5                 pkvth0dpl=0.0e-19 ku0dpl='0.50*1'            wku0dpl=7e-8                wdplku0=1 lku0dpl=11.0e-8              ldplku0=1.0                 pku0dpl=0.0e-11 keta0dpl='0.07*0'            wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0.00                wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx='0.25*1'            wku0dpx=0e-9                wdpxku0=1 lku0dpx='1.0e-8*1'          ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps='0.1*1'             wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='-0.70*1'           wku0dps=-0.0e-9             wdpsku0=1 lku0dps='9.0e-15*1'         ldpsku0=2.0                 pku0dps='-7.0e-23*0' keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps='-0.3*0'            wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa='0.01*0'            wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa='1.0e-9*0'          ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa='0.050*0'           wku0dpa=0e-7                wdpaku0=1 lku0dpa=0.0e-11             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=-0.0                wka0dpa=0                   wdpaka0=1 lka0dpa=-0.0e-7             ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa='1.5*0'             wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2='0.005*1'           wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2='3e-9*1'            ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.000               wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2='2.5e-5*1'          ldp2ku0=0.5                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2='0.5*0'             wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx='0.050*2'           wkvth0enx='8.0e-9*1'          wenxkvth0=1 lkvth0enx='1.0e-8*1'          lenxkvth0=1.0                 pkvth0enx=0 ku0enx='-0.90*1.7'         wku0enx='-0.9e-8*1.5'       wenxku0=1 lku0enx='2.0e-7*1'          lenxku0=1.0                 pku0enx='-3.0e-16*1.7' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0.0                 wka0enx=0                   wenxka0=1 lka0enx='1.0e-7*2'          lenxka0=1.0                 pka0enx='1.0e-14*1.7' kvsatenx=-0.0                wenx=0                   ku0enx0='0.15*0' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.01e-6 kvth0eny='0.04*1.7'          wkvth0eny='4.0e-10*4'         wenykvth0=1 lkvth0eny='1.0e-7*1.7'        lenykvth0=1.0                 pkvth0eny=0 ku0eny='-0.70*2'           wku0eny='-1.1e-8*1'         wenyku0=1 ku0eny0='0.025*0'           wku0eny0=0                   weny0ku0=1 lku0eny='6.0e-10*1.7'       lenyku0=1.5                 pku0eny=-0.0e-14 keta0eny=0.00                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-8             wenyka0=1 lka0eny='-6.0e-8*1.7'       lenyka0=1.0                 pka0eny='1.0e-14*1.7' kvsateny=-0.0                weny=0 kvth0eny1=0.000              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=0 ku0eny1='0.15*1.7'         wku0eny1=0.0e-8             weny1ku0=1 lku0eny1='1.0e-5*1.0'       leny1ku0=1.0                pku0eny1=-0.0e-14 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1.0                pka0eny1=0 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=-0.045              wkvth0rx=-0.0e-5             wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0.0e-16 ku0rx='0.3'               wku0rx=0.0e-8              wrxku0=1.0 lku0rx='-3.5e-10*0'        lrxku0=1                   pku0rx=0.0e-15 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.0                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=0.9027e-5           ringymin=0.117e-6 kvth0ry='-0.03*1'           wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry=0.0e-8              lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry='-0.02*1'           wku0ry=-0.0e-8             wryku0=1.0 lku0ry='-1.0e-8*1'         lryku0=1.0                 pku0ry=-0.0e-16 keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry=0                   wry=0 kvth0ry0=0.01                ku0ry0=0.02 sfxref=9.0e-8            sfxmax=3.906e-6           minwodx=0.0e-6 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0009            lkvth0odx1b=0.0e-7            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.0028           lku0odx1b=0.8e-10           lodx1bku0=1.0 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6              sfymax=10e-6             minwody=0.9e-6 wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-1.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.000            lkvth0odyb=0.0e-10           lodybkvth0=1.0 wkvth0odyb=-2.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.03             lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-1.0e-7           wodybku0=1.0               pku0odyb=0 web_mac=0  wec_mac=0 kvsatwe=0.0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_hia_mac.1 nmos ( level=54                         lmin=0.09e-06                   lmax=0.13601e-6 wmin=13.5e-06                   wmax=54.01e-06 jtsswgs='4.52e-005*(1+1.57*iboffn_flag_hia)'                               jtsswgd='4.52e-005*(1+1.57*iboffn_flag_hia)' lmin_flag=0                          lmax_flag=0                          wmin_flag=0 wmax_flag=0 tmimodel=1 )
.param ccoflag_hvt=0 rgflag_hvt=0 sigma_factor_hvt=1 rcoflag_hvt=0 scale_mos_hvt=0.9 bidirectionflag_mos_hvt=1 designflag_mos_hvt=0 iboffn_flag_hvt=0 iboffp_flag_hvt=0 totalflag_mos_hvt=1 globalflag_mos_hvt=1 mismatchflag_mos_hvt=1 global_factor_hvt=1 local_factor_hvt=1 noiseflagn_hvt=0 noiseflagp_hvt=0 noiseflagn_hvt_mc=0 noiseflagp_hvt_mc=0 sigma_factor_flicker_hvt=1
.param toxn_hvt=2.01e-009                ntoxn_hvt=1                        dxln_hvt=0 dxwn_hvt=0                        cjn_hvt=0.001686                 cjswn_hvt=1.31e-10 cjswgn_hvt=4.36e-10                 cgon_hvt=6.81825e-11              cgln_hvt=2.91624e-11 ddlcn_hvt='5.69006e-09-(5.69006e-09)' dvthn_hvt=0                        dlvthn_hvt=0 dwvthn_hvt=0                        dpvthn_hvt=0                        du0n_hvt=0 dlu0n_hvt=0                        dwu0n_hvt=0                        dpu0n_hvt=0 dvsatn_hvt=0                        dlvsatn_hvt=0                        dwvsatn_hvt=0 dpvsatn_hvt=0                        dvoffn_hvt=0                        dlvoffn_hvt=0 dwvoffn_hvt=0                        dpvoffn_hvt=0                        dagsn_hvt=0 dlagsn_hvt=0                        dwagsn_hvt=0                        dpagsn_hvt=0 dnfactorn_hvt=0                        dlnfactorn_hvt=0                        dwnfactorn_hvt=0 dpnfactorn_hvt=0                        dcitn_hvt=0                        dlcitn_hvt=0 dwcitn_hvt=0                        dpcitn_hvt=0                        deta0n_hvt=0 dleta0n_hvt=0                        dweta0n_hvt=0                        dpeta0n_hvt=0 dk2n_hvt=0                        dlk2n_hvt=0                        dpclmn_hvt=0 dlpclmn_hvt=0                        dwpclmn_hvt=0                        dppclmn_hvt=0 dua1n_hvt=0                        dlua1n_hvt=0                        dwua1n_hvt=0 dpua1n_hvt=0                        datn_hvt=0                        dlatn_hvt=0 dwatn_hvt=0                        dpatn_hvt=0                        dkt1n_hvt=0 dlkt1n_hvt=0                        dwkt1n_hvt=0                        dpkt1n_hvt=0 dkt2n_hvt=0                        duc1n_hvt=0                        cfn_hvt='6.62e-11+9.73e-11*ccoflag_hvt' jtsswgn_hvt='7.6e-006*(1+0.645*iboffn_flag_hvt)' dpdiblc2n_hvt=0                        dminvn_hvt=0 da0n_hvt=0 ss_flagn_hvt=0 ff_flagn_hvt=0 sf_flagn_hvt=0 fs_flagn_hvt=0
.param toxp_hvt=2.18e-009                ntoxp_hvt=1                        dxlp_hvt=0 dxwp_hvt=0                        cjp_hvt=0.001739                 cjswp_hvt=1.242e-10 cjswgp_hvt=3e-10                    cgop_hvt=4.92779e-11              cglp_hvt=4.63343e-11 ddlcp_hvt='5.66905e-09-(5.66905e-09)' dvthp_hvt=0                        dlvthp_hvt=0 dwvthp_hvt=0                        dpvthp_hvt=0                        dk2p_hvt=0 dlk2p_hvt=0                        dwk2p_hvt=0                        dpk2p_hvt=0 deta0p_hvt=0                        dleta0p_hvt=0                        dweta0p_hvt=0 dpeta0p_hvt=0                        dvoffp_hvt=0                        dlvoffp_hvt=0 dwvoffp_hvt=0                        dpvoffp_hvt=0                        dcitp_hvt=0 dlcitp_hvt=0                        dwcitp_hvt=0                        dpcitp_hvt=0 dnfactorp_hvt=0                        dlnfactorp_hvt=0                        dwnfactorp_hvt=0 dpnfactorp_hvt=0                        du0p_hvt=0                        dlu0p_hvt=0 dwu0p_hvt=0                        dpu0p_hvt=0                        dubp_hvt=0 dlubp_hvt=0                        dwubp_hvt=0                        dpubp_hvt=0 dpclmp_hvt=0                        dlpclmp_hvt=0                        dwpclmp_hvt=0 dppclmp_hvt=0                        dvsatp_hvt=0                        dlvsatp_hvt=0 dwvsatp_hvt=0                        dpvsatp_hvt=0                        da0p_hvt=0 dla0p_hvt=0                        dwa0p_hvt=0                        dpa0p_hvt=0 dagsp_hvt=0                        dlagsp_hvt=0                        dwagsp_hvt=0 dpagsp_hvt=0                        dpkt1p_hvt=0                        datp_hvt=0 dlatp_hvt=0                        dwatp_hvt=0                        dpatp_hvt=0 dua1p_hvt=0                        dlua1p_hvt=0                        dwua1p_hvt=0 dpua1p_hvt=0                        cfp_hvt='9e-11+0.92e-10*ccoflag_hvt' jtsswgp_hvt='4.5e-007*(1+0.42*iboffp_flag_hvt)' dpdiblc2p_hvt=0                        dminvp_hvt=0 dketap_hvt=0                        dlketap_hvt=0                        dwketap_hvt=0 dpketap_hvt=0 ss_flagp_hvt=0 ff_flagp_hvt=0 sf_flagp_hvt=0 fs_flagp_hvt=0 monte_flagn_hvt=0 monte_flagp_hvt=0 c1fn_hvt=1.57e+042                c2fn_hvt=3.13e+025                c3fn_hvt=2.21e+009 c1fp_hvt=2.66e+042                c2fp_hvt=8.23e+026                c3fp_hvt=2.03e+010
.param ccoflag_lvt=0 rgflag_lvt=0 sigma_factor_lvt=1 rcoflag_lvt=0 scale_mos_lvt=0.9 bidirectionflag_mos_lvt=1 designflag_mos_lvt=0 iboffn_flag_lvt=0 totalflag_mos_lvt=1 globalflag_mos_lvt=1 mismatchflag_mos_lvt=1 global_factor_lvt=1 local_factor_lvt=1 iboffp_flag_lvt=0 noiseflagn_lvt=0 noiseflagp_lvt=0 noiseflagn_lvt_mc=0 noiseflagp_lvt_mc=0 sigma_factor_flicker_lvt=1
.param toxn_lvt=1.95e-009                dxln_lvt=0                        dxwn_lvt=0 cjn_lvt=0.00139                  cjswn_lvt=1.050e-10                cjswgn_lvt=2.890e-10 cgon_lvt=9.775e-011               cgln_lvt=1.449e-011               ddlcn_lvt='6.25e-009-(6.25e-009)' ntoxn_lvt=1                        cfn_lvt='6.62e-011+9.73e-11*ccoflag_lvt' dvthn_lvt=0                        dlvthn_lvt=0                        dwvthn_lvt=0 dpvthn_lvt=0                        du0n_lvt=0                        dlu0n_lvt=0 dwu0n_lvt=0                        dpu0n_lvt=0                        dvsatn_lvt=0 dlvsatn_lvt=0                        dwvsatn_lvt=0                        dpvsatn_lvt=0 dk2n_lvt=0                        dlk2n_lvt=0                        dwk2n_lvt=0 dpk2n_lvt=0                        dvoffn_lvt=0                        dlvoffn_lvt=0 dwvoffn_lvt=0                        dpvoffn_lvt=0                        dpdiblc2n_lvt=0 dlpdiblc2n_lvt=0                        dwpdiblc2n_lvt=0                        dppdiblc2n_lvt=0 dagsn_lvt=0                        dlagsn_lvt=0                        dwagsn_lvt=0 dpagsn_lvt=0                        deta0n_lvt=0                        dleta0n_lvt=0 dweta0n_lvt=0                        dpeta0n_lvt=0                        dpclmn_lvt=0 dlpclmn_lvt=0                        dwpclmn_lvt=0                        dppclmn_lvt=0 dminvn_lvt=0                        dua1n_lvt=0                        datn_lvt=0 dlatn_lvt=0                        dwatn_lvt=0                        dpatn_lvt=0 jtsswgn_lvt='5.2e-006*(1+1.55*iboffn_flag_lvt)' ss_flagn_lvt=0 ff_flagn_lvt=0 sf_flagn_lvt=0 fs_flagn_lvt=0 monte_flagn_lvt=0
.param toxp_lvt=2.18e-009                dxlp_lvt=0                        dxwp_lvt=0 cgop_lvt=5.71e-011                cglp_lvt=6.7e-011                 ddlcp_lvt='7.64e-009-(7.64e-009)' cjp_lvt=0.001474                 cjswp_lvt=1.070e-10                cjswgp_lvt=2.070e-10 cfp_lvt='9e-011+9.2e-11*ccoflag_lvt' dvthp_lvt=0 dlvthp_lvt=0                        dwvthp_lvt=0                        dpvthp_lvt=0 dk2p_lvt=0                        dlk2p_lvt=0                        dwk2p_lvt=0 dpk2p_lvt=0                        deta0p_lvt=0                        dweta0p_lvt=0 dvoffp_lvt=0                        dlvoffp_lvt=0                        dwvoffp_lvt=0 dpvoffp_lvt=0                        du0p_lvt=0                        dlu0p_lvt=0 dwu0p_lvt=0                        dpu0p_lvt=0                        dpclmp_lvt=0 dlpclmp_lvt=0                        dwpclmp_lvt=0                        dppclmp_lvt=0 dpdiblc2p_lvt=0                        dwpdiblc2p_lvt=0                        dlpdiblc2p_lvt=0 dppdiblc2p_lvt=0                        da0p_lvt=0                        dla0p_lvt=0 dwa0p_lvt=0                        dpa0p_lvt=0                        dagsp_lvt=0 dlagsp_lvt=0                        dwagsp_lvt=0                        dpagsp_lvt=0 ntoxp_lvt=1                        dvsatp_lvt=0                        dlvsatp_lvt=0 dwvsatp_lvt=0                        dpvsatp_lvt=0                        dminvp_lvt=0 datp_lvt=0                        dua1p_lvt=0                        dlua1p_lvt=0 dwua1p_lvt=0                        dpua1p_lvt=0 jtsswgp_lvt='7.8e-006*(1+0.3*iboffp_flag_lvt)' ss_flagp_lvt=0 ff_flagp_lvt=0 sf_flagp_lvt=0 fs_flagp_lvt=0 monte_flagp_lvt=0 c1fn_lvt=8.20e+041                c2fn_lvt=7.70e+023                c3fn_lvt=4.57e+006 c1fp_lvt=2.03e+042                c2fp_lvt=3.23e+026                c3fp_lvt=2.00e+010
.param scale_cap=0.9 ccoflag_cap=0
.param cgminn_var=1       dcgn_var=1           cfrwn_var=1           cfrln_var=1 dvgsn_var_a=1     dvgsn_var_w=0       dvgsn_var_l=0 dxln_var=0         dxwn_var=0 x_facn_var=0
.param cgminp_var=1                 dcgp_var=1                 cfrwp_var=1                 cfrlp_var=1 dvgsp_var_a=1                 dvgsp_var_w=0                 dvgsp_var_l=0 dxlp_var=0                 dxwp_var=0 x_facp_var=0
.subckt nmoscap ng nds lr=1u wr=1u scale=scale_cap _ccoflag_cap=ccoflag_cap multi=1
.param xl_mvar=4.785e-09
.param xw_mvar=-3.464e-08
.param area_mvar='(lr*scale-xl_mvar+dxln_var)*(wr*scale-xw_mvar+dxwn_var)'
.param cf_mvar='(3.10e-11+9.73e-11*_ccoflag_cap)*cfrwn_var*2*(wr*scale-xw_mvar+dxwn_var)+(9.525e-11)*cfrln_var*2*(lr*scale-xl_mvar+dxln_var)'
.param cgmin_mvar='(2.661e-03)*cgminn_var*(1+(-3.531e-04)*(temper-25))*area_mvar'
.param dcg_mvar='(1.582e-02)*(1+(0.000e+00)/(wr*scale-xw_mvar+dxwn_var)+(0.000e+00)/(lr*scale-xl_mvar+dxln_var)+(0.000e+00)/(area_mvar))*dcgn_var*area_mvar'
.param dvgs1_mvar='dvgsn_var_a+dvgsn_var_w*1e-6/(wr*scale-xw_mvar+dxwn_var)+dvgsn_var_l*1e-6/(lr*scale-xl_mvar+dxln_var)'
.param dvgs_mvar='-0.0549*(1+(3.664e-03)*(temper-25))*dvgs1_mvar'
.param vgnorm_mvar='2.533e-03*(1+(7.475e-03)*(temper-25))'
.param delta1_mvar=0.26279
.param delta2_mvar=0.26404
.param dis1_mvar=1.18267
.param dis2_mvar=0.02154
cg ng nds 'multi*(cf_mvar+cgmin_mvar+dcg_mvar*(0.5+(vgnorm_mvar*(pwr((v(ng,nds)-(dvgs_mvar-dis1_mvar))*(v(ng,nds)-(dvgs_mvar-dis1_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis1_mvar))*(v(ng,nds)-(dvgs_mvar+dis1_mvar))+delta1_mvar*delta1_mvar,0.5))+pwr((v(ng,nds)-(dvgs_mvar-dis2_mvar))*(v(ng,nds)-(dvgs_mvar-dis2_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis2_mvar))*(v(ng,nds)-(dvgs_mvar+dis2_mvar))+delta2_mvar*delta2_mvar,0.5))/(4*(dis2_mvar+vgnorm_mvar*dis1_mvar))))'
.param for_eff_mvar='2.625e+04*pwr(abs((273.15+temper)/(273.15+25)),0.531)'
.param varbf_mvar=8.292
.param rev_eff_mvar='2.642e+04*pwr(abs((273.15+temper)/(273.15+25)),0.451)'
.param varbr_mvar=1.875
.param a1_mvar=1.766
.param a2_mvar=426.995
.param a3_mvar='-187613.139*pwr(abs((273.15+temper)/(273.15+25)),0.431)'
.param a_mvar=1.012
.param area1_mvar='(lr*scale-xl_mvar+dxln_var)*(pwr(abs(wr*scale*1e6-xw_mvar*1e6+dxwn_var*1e6),a_mvar))*1e-6'
gdf1 ng nds cur='multi*(exp(x_facn_var)*area1_mvar*(for_eff_mvar*(pwr(0.5*(sqrt(v(ng,nds)*v(ng,nds)+a1_mvar)+v(ng,nds)),varbf_mvar)-pwr(abs(0.5*pwr(abs(a1_mvar),0.5)),varbf_mvar))-rev_eff_mvar*(pwr(0.5*(sqrt(v(ng,nds)*v(ng,nds)+a2_mvar)-v(ng,nds)),varbr_mvar)-pwr(abs(0.5*pwr(abs(a2_mvar),0.5)),varbr_mvar))+a3_mvar*v(ng,nds)))'
.ends nmoscap
.subckt pmoscap ng nds lr=1u wr=1u scale=scale_cap _ccoflag_cap=ccoflag_cap multi=1
.param xl_mvar=1.227e-08
.param xw_mvar=-4.074e-08
.param area_mvar='(lr*scale-xl_mvar+dxlp_var)*(wr*scale-xw_mvar+dxwp_var)'
.param cf_mvar='(6.409e-12+0.92e-10*_ccoflag_cap)*cfrwp_var*2*(wr*scale-xw_mvar+dxwp_var)+(1.493e-21)*cfrlp_var*2*(lr*scale-xl_mvar+dxlp_var)'
.param cgmin_mvar='(2.300e-03)*cgminp_var*(1+(2.0e-04)*(temper-25))*area_mvar'
.param dcg_mvar='(1.309e-02)*(1+(0.000e+00)/(wr*scale-xw_mvar+dxwp_var)+(0.000e+00)/(lr*scale-xl_mvar+dxlp_var)+(0.000e+00)/(area_mvar))*dcgp_var*area_mvar'
.param dvgs1_mvar='dvgsp_var_a+dvgsp_var_w*1e-6/(wr*scale-xw_mvar+dxwp_var)+dvgsp_var_l*1e-6/(lr*scale-xl_mvar+dxlp_var)'
.param dvgs_mvar='0.1244*(1+(2.845e-03)*(temper-25))*dvgs1_mvar'
.param vgnorm_mvar='1.606e-02*(1+(6.809e-03)*(temper-25))'
.param delta1_mvar=0.248866
.param delta2_mvar=0.248857
.param dis1_mvar=0.525249
.param dis2_mvar=0.007000
cg ng nds 'multi*(cf_mvar+cgmin_mvar+dcg_mvar*(0.5-(vgnorm_mvar*(pwr((v(ng,nds)-(dvgs_mvar-dis1_mvar))*(v(ng,nds)-(dvgs_mvar-dis1_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis1_mvar))*(v(ng,nds)-(dvgs_mvar+dis1_mvar))+delta1_mvar*delta1_mvar,0.5))+pwr((v(ng,nds)-(dvgs_mvar-dis2_mvar))*(v(ng,nds)-(dvgs_mvar-dis2_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis2_mvar))*(v(ng,nds)-(dvgs_mvar+dis2_mvar))+delta2_mvar*delta2_mvar,0.5))/(4*(dis2_mvar+vgnorm_mvar*dis1_mvar))))'
.param for_eff_mvar='1.321e+04*pwr(abs((273.15+temper)/(273.15+25)),0.538)'
.param varbf_mvar=5.315
.param rev_eff_mvar='2.671e+04*pwr(abs((273.15+temper)/(273.15+25)),0.478)'
.param varbr_mvar=1.000
.param a1_mvar=0.176
.param a2_mvar=2.025
.param a3_mvar='-20540.928*pwr(abs((273.15+temper)/(273.15+25)),0.447)'
.param a_mvar=1.027
.param area1_mvar='(lr*scale-xl_mvar+dxlp_var)*(pwr(abs(wr*scale*1e6-xw_mvar*1e6+dxwp_var*1e6),a_mvar))*1e-6'
gdf1 ng nds cur='multi*(exp(x_facp_var)*area1_mvar*(rev_eff_mvar*(pwr(0.5*(sqrt(v(ng,nds)*v(ng,nds)+a1_mvar)+v(ng,nds)),varbr_mvar)-pwr(abs(0.5*pwr(abs(a1_mvar),0.5)),varbr_mvar))-for_eff_mvar*(pwr(0.5*(sqrt(v(ng,nds)*v(ng,nds)+a2_mvar)-v(ng,nds)),varbf_mvar)-pwr(abs(0.5*pwr(abs(a2_mvar),0.5)),varbf_mvar))+a3_mvar*v(ng,nds)))'
.ends pmoscap
.param scale_cap_12=0.9 ccoflag_cap_12=0
.param cgminn_var12=1       dcgn_var12=1           cfrwn_var12=1           cfrln_var12=1 dvgsn_var12_a=1     dvgsn_var12_w=0       dvgsn_var12_l=0 dxln_var12=0         dxwn_var12=0 x_facn_var12=0
.subckt nmoscap_12 ng nds lr=1u wr=1u scale=scale_cap_12 _ccoflag_cap=ccoflag_cap_12 multi=1
.param xl_mvar=8.269e-09
.param xw_mvar=-4.075e-08
.param area_mvar='(lr*scale-xl_mvar+dxln_var12)*(wr*scale-xw_mvar+dxwn_var12)'
.param cf_mvar='(2.8e-11+9.3e-11*_ccoflag_cap)*cfrwn_var12*2*(wr*scale-xw_mvar+dxwn_var12)+(7.379e-11)*cfrln_var12*2*(lr*scale-xl_mvar+dxln_var12)'
.param cgmin_mvar='(2.442e-03)*cgminn_var12*(1+(1.921e-04)*(temper-25))*area_mvar'
.param dcg_mvar='(1.222e-02)*(1+(0.000e+00)/(wr*scale-xw_mvar+dxwn_var12)+(0.000e+00)/(lr*scale-xl_mvar+dxln_var12)+(0.000e+00)/(area_mvar))*dcgn_var12*area_mvar'
.param dvgs1_mvar='dvgsn_var12_a+dvgsn_var12_w*1e-6/(wr*scale-xw_mvar+dxwn_var12)+dvgsn_var12_l*1e-6/(lr*scale-xl_mvar+dxln_var12)'
.param dvgs_mvar='-0.0762*(1+(2.023e-03)*(temper-25))*dvgs1_mvar'
.param vgnorm_mvar='-9.463e-02*(1+(-1.288e-03)*(temper-25))'
.param delta1_mvar=0.44631
.param delta2_mvar=0.44577
.param dis1_mvar=0.22284
.param dis2_mvar=0.03146
cg ng nds 'multi*(cf_mvar+cgmin_mvar+dcg_mvar*(0.5+(vgnorm_mvar*(pwr((v(ng,nds)-(dvgs_mvar-dis1_mvar))*(v(ng,nds)-(dvgs_mvar-dis1_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis1_mvar))*(v(ng,nds)-(dvgs_mvar+dis1_mvar))+delta1_mvar*delta1_mvar,0.5))+pwr((v(ng,nds)-(dvgs_mvar-dis2_mvar))*(v(ng,nds)-(dvgs_mvar-dis2_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis2_mvar))*(v(ng,nds)-(dvgs_mvar+dis2_mvar))+delta2_mvar*delta2_mvar,0.5))/(4*(dis2_mvar+vgnorm_mvar*dis1_mvar))))'
.param for_eff_mvar='4.962e+02*pwr(abs((273.15+temper)/(273.15+25)),0.724)'
.param varbf_mvar=4.939
.param rev_eff_mvar='7.450e+01*pwr(abs((273.15+temper)/(273.15+25)),0.523)'
.param varbr_mvar=2.030
.param a1_mvar=0.273
.param a2_mvar=38.942
.param a3_mvar='-242.495*pwr(abs((273.15+temper)/(273.15+25)),0.497)'
.param a_mvar=0.945
.param area1_mvar='(lr*scale-xl_mvar+dxln_var12)*(pwr(abs(wr*scale*1e6-xw_mvar*1e6+dxwn_var12*1e6),a_mvar))*1e-6'
gdf1 ng nds cur='multi*(exp(x_facn_var12)*area1_mvar*(for_eff_mvar*(pwr(0.5*(sqrt(v(ng,nds)*v(ng,nds)+a1_mvar)+v(ng,nds)),varbf_mvar)-pwr(abs(0.5*pwr(abs(a1_mvar),0.5)),varbf_mvar))-rev_eff_mvar*(pwr(0.5*(sqrt(v(ng,nds)*v(ng,nds)+a2_mvar)-v(ng,nds)),varbr_mvar)-pwr(abs(0.5*pwr(abs(a2_mvar),0.5)),varbr_mvar))+a3_mvar*v(ng,nds)))'
.ends nmoscap_12
.param scale_cap_18=0.9 ccoflag_cap_18=0
.param cgminn_var18=1       dcgn_var18=1           cfrwn_var18=1           cfrln_var18=1 dvgsn_var18_a=1     dvgsn_var18_w=0       dvgsn_var18_l=0 dxln_var18=0         dxwn_var18=0
.param cgminp_var18=1                 dcgp_var18=1                 cfrwp_var18=1                 cfrlp_var18=1 dvgsp_var18_a=1                 dvgsp_var18_w=0                 dvgsp_var18_l=0 dxlp_var18=0                 dxwp_var18=0
.subckt nmoscap_18 ng nds lr=1u wr=1u scale=scale_cap_18 _ccoflag_cap=ccoflag_cap_18 multi=1
.param xl_mvar=-4.832e-09
.param xw_mvar=-3.917e-08
.param area_mvar='(lr*scale-xl_mvar+dxln_var18)*(wr*scale-xw_mvar+dxwn_var18)'
.param cf_mvar='(6.978e-11+5.742e-11*_ccoflag_cap)*cfrwn_var18*2*(wr*scale-xw_mvar+dxwn_var18)+(9.066e-11)*cfrln_var18*2*(lr*scale-xl_mvar+dxln_var18)'
.param cgmin_mvar='(1.516e-03)*cgminn_var18*(1+(0.000e+00)*(temper-25))*area_mvar'
.param dcg_mvar='(8.784e-03)*(1+(0.000e+00)/(wr*scale-xw_mvar+dxwn_var18)+(0.000e+00)/(lr*scale-xl_mvar+dxln_var18)+(0.000e+00)/(area_mvar))*dcgn_var18*area_mvar'
.param dvgs1_mvar='dvgsn_var18_a+dvgsn_var18_w*1e-6/(wr*scale-xw_mvar+dxwn_var18)+dvgsn_var18_l*1e-6/(lr*scale-xl_mvar+dxln_var18)'
.param dvgs_mvar='-0.0647*(1+(0.000e+00)*(temper-25))*dvgs1_mvar'
.param vgnorm_mvar='-2.096e+00*(1+(0.000e+00)*(temper-25))'
.param delta1_mvar=0.36109
.param delta2_mvar=0.35891
.param dis1_mvar=-0.018
.param dis2_mvar=0.019
cg ng nds 'multi*(cf_mvar+cgmin_mvar+dcg_mvar*(0.5+(vgnorm_mvar*(pwr((v(ng,nds)-(dvgs_mvar-dis1_mvar))*(v(ng,nds)-(dvgs_mvar-dis1_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis1_mvar))*(v(ng,nds)-(dvgs_mvar+dis1_mvar))+delta1_mvar*delta1_mvar,0.5))+pwr((v(ng,nds)-(dvgs_mvar-dis2_mvar))*(v(ng,nds)-(dvgs_mvar-dis2_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis2_mvar))*(v(ng,nds)-(dvgs_mvar+dis2_mvar))+delta2_mvar*delta2_mvar,0.5))/(4*(dis2_mvar+vgnorm_mvar*dis1_mvar))))'
.ends nmoscap_18
.subckt pmoscap_18 ng nds lr=1u wr=1u scale=scale_cap_18 _ccoflag_cap=ccoflag_cap_18 multi=1
.param xl_mvar=-4.530e-09
.param xw_mvar=-5.150e-08
.param area_mvar='(lr*scale-xl_mvar+dxlp_var18)*(wr*scale-xw_mvar+dxwp_var18)'
.param cf_mvar='(4.357e-22+5.68e-11*_ccoflag_cap)*cfrwp_var18*2*(wr*scale-xw_mvar+dxwp_var18)+(2.453e-21)*cfrlp_var18*2*(lr*scale-xl_mvar+dxlp_var18)'
.param cgmin_mvar='(1.280e-03)*cgminp_var18*(1+(0)*(temper-25))*area_mvar'
.param dcg_mvar='(7.932e-03)*(1+(0.000e+00)/(wr*scale-xw_mvar+dxwp_var18)+(0.000e+00)/(lr*scale-xl_mvar+dxlp_var18)+(0.000e+00)/(area_mvar))*dcgp_var18*area_mvar'
.param dvgs1_mvar='dvgsp_var18_a+dvgsp_var18_w*1e-6/(wr*scale-xw_mvar+dxwp_var18)+dvgsp_var18_l*1e-6/(lr*scale-xl_mvar+dxlp_var18)'
.param dvgs_mvar='0.2781*(1+(0)*(temper-25))*dvgs1_mvar'
.param vgnorm_mvar='5.762e-03*(1+(0)*(temper-25))'
.param delta1_mvar=0.322108
.param delta2_mvar=0.322500
.param dis1_mvar=0.804810
.param dis2_mvar=0.007000
cg ng nds 'multi*(cf_mvar+cgmin_mvar+dcg_mvar*(0.5-(vgnorm_mvar*(pwr((v(ng,nds)-(dvgs_mvar-dis1_mvar))*(v(ng,nds)-(dvgs_mvar-dis1_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis1_mvar))*(v(ng,nds)-(dvgs_mvar+dis1_mvar))+delta1_mvar*delta1_mvar,0.5))+pwr((v(ng,nds)-(dvgs_mvar-dis2_mvar))*(v(ng,nds)-(dvgs_mvar-dis2_mvar))+delta1_mvar*delta1_mvar,0.5)-pwr((v(ng,nds)-(dvgs_mvar+dis2_mvar))*(v(ng,nds)-(dvgs_mvar+dis2_mvar))+delta2_mvar*delta2_mvar,0.5))/(4*(dis2_mvar+vgnorm_mvar*dis1_mvar))))'
.ends pmoscap_18
.param ccoflag_na=0 rgflag_na=0 rcoflag_na=0 scale_mos_na=0.9 sigma_factor_na=1 totalflag_mos_na=1 globalflag_mos_na=1 mismatchflag_mos_na=1 global_factor_na=1 local_factor_na=1 noiseflagn_na=0 noiseflagn_na_mc=0 sigma_factor_flicker_na=1
.param toxn_na=1.96e-009                dxln_na=0                        dxwn_na=0 cjn_na=0.000159                 cjswn_na=1.99e-010                cjswgn_na=1.49e-010 cgon_na=8.8e-011                 cgln_na=3.0012e-010              ddlcn_na='1.94e-008-(1.94e-008)' cfn_na='6.22e-011+9.73e-11*ccoflag_na' dvthn_na=0                        dlvthn_na=0 dwvthn_na=0                        dpvthn_na=0                        du0n_na=0 dlu0n_na=0                        dwu0n_na=0                        dpu0n_na=0 dlk2n_na=0                        dwk2n_na=0                        dpk2n_na=0 dvsatn_na=0                        dlvsatn_na=0                        dwvsatn_na=0 dpvsatn_na=0                        dpdiblc2n_na=0                        dlpdiblc2n_na=0 dwpdiblc2n_na=0                        dppdiblc2n_na=0                        ntoxn_na=1 dagsn_na=0                        dlagsn_na=0                        dwagsn_na=0 dpagsn_na=0                        dua1n_na=0 monte_flagn_na=0 c1fn_na=9e+041                   c2fn_na=5.65e+022                c3fn_na=8.53e+06
.param ccoflag_na12=0 sigma_factor_na12=1 rgflag_na12=0 rcoflag_na12=0 scale_mos_na12=0.9 totalflag_mos_na12=1 globalflag_mos_na12=1 mismatchflag_mos_na12=1 global_factor_na12=1 local_factor_na12=1 noiseflagn_na12=0 noiseflagn_na12_mc=0 sigma_factor_flicker_na12=1
.param toxn_na12=2.43e-09                 dxln_na12=0                        dxwn_na12=0 cgon_na12=1.7433e-010              cgln_na12=4e-011                   ddlcn_na12='1.2924e-08-(1.2924e-08)' cjn_na12=0.0001576                cjswn_na12=2.102e-10                cjswgn_na12=1.551e-10 cfn_na12='6.7e-11+9.3e-11*ccoflag_na12' dvthn_na12=0 dlvthn_na12=0                        dwvthn_na12=0                        dpvthn_na12=0 du0n_na12=0                        dlu0n_na12=0                        dwu0n_na12=0 dpu0n_na12=0                        dvsatn_na12=0                        dwvsatn_na12=0 dk2n_na12=0                        dlk2n_na12=0                        dwk2n_na12=0 dpk2n_na12=0                        deta0n_na12=0                        dweta0n_na12=0 dagsn_na12=0                        dlagsn_na12=0                        dwagsn_na12=0 dpagsn_na12=0                        dvoffn_na12=0                        dlvoffn_na12=0 dwvoffn_na12=0                        dpvoffn_na12=0                        dcitn_na12=0 dlcitn_na12=0                        dwcitn_na12=0                        dpcitn_na12=0 duan_na12=0                        dluan_na12=0                        dwuan_na12=0 dpuan_na12=0                        dubn_na12=0                        dlubn_na12=0 dwubn_na12=0                        dpubn_na12=0                        dkt1n_na12=0 dlkt1n_na12=0                        dwkt1n_na12=0                        dpkt1n_na12=0 datn_na12=0                        dlatn_na12=0                        dwatn_na12=0 dpatn_na12=0                        dpdiblc2n_na12=0                        dlpdiblc2n_na12=0 dwpdiblc2n_na12=0                        dppdiblc2n_na12=0                        dlvsatn_na12=0 dpvsatn_na12=0                        da0n_na12=0                        dla0n_na12=0 dwa0n_na12=0                        dpa0n_na12=0 ntoxn_na12=1                        dpclmn_na12=0                        dlpclmn_na12=0 dwpclmn_na12=0                        dppclmn_na12=0                        duc1n_na12=0 dluc1n_na12=0                        dwuc1n_na12=0                        dpuc1n_na12=0 ff_flagn_na12=0 monte_flagn_na12=0 c1fn_na12=3.00000e+42              c2fn_na12=4.330000e+22             c3fn_na12=1.120000e+06
.param ccoflag_na18=0 sigma_factor_na18=1 rcoflag_na18=0 scale_mos_na18=0.9 rgflag_na18=0 totalflag_mos_na18=1 globalflag_mos_na18=1 mismatchflag_mos_na18=1 global_factor_na18=1 local_factor_na18=1 noiseflagn_na18=0 noiseflagn_na18_mc=0 sigma_factor_flicker_na18=1
.param toxn_na18=3.36e-09                 dxln_na18=0                        dxwn_na18=0 cjn_na18=0.000161                 cjswn_na18=2.08e-10                 cjswgn_na18=1.62e-10 cgon_na18=4.925043e-11             cgln_na18=3.247859e-10             ddlcn_na18='3.542614e-08-(3.542614e-08)' dvthn_na18=0                        dlvthn_na18=0                        dwvthn_na18=0 dpvthn_na18=0                        cfn_na18='8.050e-11+7.81e-11*ccoflag_na18' du0n_na18=0                        dlu0n_na18=0                        dwu0n_na18=0 dpu0n_na18=0                        dvsatn_na18=0                        dlvsatn_na18=0 dwvsatn_na18=0                        dpvsatn_na18=0                        dk2n_na18=0 drdswn_na18=0                        dvoffn_na18=0                        dlvoffn_na18=0 dwvoffn_na18=0                        dpvoffn_na18=0                        dpdiblc2n_na18=0 dlpdiblc2n_na18=0                        dwpdiblc2n_na18=0                        dppdiblc2n_na18=0 dagsn_na18=0                        dlagsn_na18=0                        dwagsn_na18=0 dpagsn_na18=0                        dnfactorn_na18=0                        dlnfactorn_na18=0 dwnfactorn_na18=0                        dpnfactorn_na18=0                        dcitn_na18=0 dlcitn_na18=0                        dwcitn_na18=0                        dpcitn_na18=0 deta0n_na18=0                        dleta0n_na18=0                        dweta0n_na18=0 dpeta0n_na18=0                        dub1n_na18=0                        dlk2n_na18=0 dwk2n_na18=0                        dpk2n_na18=0                        dkt1n_na18=0 dlkt2n_na18=0                        dla0n_na18=0                        dwa0n_na18=0 dlucn_na18=0                        dlketan_na18=0 monte_flagn_na18=0 c1fn_na18=8.520000e+41             c2fn_na18=3.000000e+24             c3fn_na18=9.160000e+07
.param ccoflag_na18ud15=0 sigma_factor_na18ud15=1 rcoflag_na18ud15=0 scale_mos_na18ud15=0.9 rgflag_na18ud15=0 totalflag_mos_na18ud15=1 globalflag_mos_na18ud15=1 mismatchflag_mos_na18ud15=1 global_factor_na18ud15=1 local_factor_na18ud15=1 noiseflagn_na18ud15=0 noiseflagn_na18ud15_mc=0 sigma_factor_flicker_na18ud15=1
.param toxn_na18ud15=3.36e-09                 dxln_na18ud15=0                        dxwn_na18ud15=0 cjn_na18ud15=0.000161                 cjswn_na18ud15=2.08e-10                 cjswgn_na18ud15=1.62e-10 cgon_na18ud15=4.925043e-11             cgln_na18ud15=3.247859e-10             ddlcn_na18ud15='3.542614e-08-(3.542614e-08)' dvthn_na18ud15=0                        dlvthn_na18ud15=0                        dwvthn_na18ud15=0 dpvthn_na18ud15=0                        cfn_na18ud15='8.050e-11+7.81e-11*ccoflag_na18ud15' du0n_na18ud15=0                        dlu0n_na18ud15=0                        dwu0n_na18ud15=0 dpu0n_na18ud15=0                        dvsatn_na18ud15=0                        dlvsatn_na18ud15=0 dwvsatn_na18ud15=0                        dpvsatn_na18ud15=0                        dk2n_na18ud15=0 drdswn_na18ud15=0                        dvoffn_na18ud15=0                        dlvoffn_na18ud15=0 dwvoffn_na18ud15=0                        dpvoffn_na18ud15=0                        dpdiblc2n_na18ud15=0 dlpdiblc2n_na18ud15=0                        dwpdiblc2n_na18ud15=0                        dppdiblc2n_na18ud15=0 dagsn_na18ud15=0                        dlagsn_na18ud15=0                        dwagsn_na18ud15=0 dpagsn_na18ud15=0                        dnfactorn_na18ud15=0                        dlnfactorn_na18ud15=0 dwnfactorn_na18ud15=0                        dpnfactorn_na18ud15=0                        dcitn_na18ud15=0 dlcitn_na18ud15=0                        dwcitn_na18ud15=0                        dpcitn_na18ud15=0 deta0n_na18ud15=0                        dleta0n_na18ud15=0                        dweta0n_na18ud15=0 dpeta0n_na18ud15=0                        dub1n_na18ud15=0                        dlk2n_na18ud15=0 dwk2n_na18ud15=0                        dpk2n_na18ud15=0                        dkt1n_na18ud15=0 dlkt2n_na18ud15=0                        dla0n_na18ud15=0                        dwa0n_na18ud15=0 dlucn_na18ud15=0                        dlketan_na18ud15=0 monte_flagn_na18ud15=0 c1fn_na18ud15=8.520000e+41             c2fn_na18ud15=3.000000e+24             c3fn_na18ud15=9.160000e+07
.param toxn_ms_global=0 dxln_ms_global=0 dxwn_ms_global=0 cjn_ms_global=0 cjswn_ms_global=0 cjswgn_ms_global=0 cgon_ms_global=0 cgln_ms_global=0 cfn_ms_global=0 ntoxn_ms_global=0 dvthn_ms_global=0 dlvthn_ms_global=0 dwvthn_ms_global=0 dpvthn_ms_global=0 du0n_ms_global=0 dlu0n_ms_global=0 dwu0n_ms_global=0 dpu0n_ms_global=0 dvsatn_ms_global=0 dlvsatn_ms_global=0 dwvsatn_ms_global=0 dpvsatn_ms_global=0 dk2n_ms_global=0 dlk2n_ms_global=0 dwk2n_ms_global=0 dlvoffn_ms_global=0 dpvoffn_ms_global=0 dpdiblc2n_ms_global=0 dppdiblc2n_ms_global=0 dagsn_ms_global=0 dwagsn_ms_global=0 dlcitn_ms_global=0 dpcitn_ms_global=0 dpclmn_ms_global=0 dminvn_ms_global=0 dketan_ms_global=0 dlketan_ms_global=0 dpketan_ms_global=0 dua1n_ms_global=0 datn_ms_global=0 ss_flagn_ms_global=0 ff_flagn_ms_global=0 monte_flagn_ms_global=0 deta0n_ms_global=0 sf_flagn_ms_global=0 fs_flagn_ms_global=0 toxp_ms_global=0 dxlp_ms_global=0 dxwp_ms_global=0 cjp_ms_global=0 cjswp_ms_global=0 cjswgp_ms_global=0 cgop_ms_global=0 cglp_ms_global=0 cfp_ms_global=0 ntoxp_ms_global=0 dvthp_ms_global=0 dlvthp_ms_global=0 dwvthp_ms_global=0 dpvthp_ms_global=0 dk2p_ms_global=0 dlk2p_ms_global=0 deta0p_ms_global=0 dlvoffp_ms_global=0 dpvoffp_ms_global=0 du0p_ms_global=0 dlu0p_ms_global=0 dwu0p_ms_global=0 dpu0p_ms_global=0 dlpclmp_ms_global=0 dpdiblc2p_ms_global=0 dvsatp_ms_global=0 dlvsatp_ms_global=0 dwvsatp_ms_global=0 dpvsatp_ms_global=0 dagsp_ms_global=0 dwagsp_ms_global=0 dminvp_ms_global=0 datp_ms_global=0 dpatp_ms_global=0 dua1p_ms_global=0 dpua1p_ms_global=0 dketap_ms_global=0 dpketap_ms_global=0 ss_flagp_ms_global=0 ff_flagp_ms_global=0 monte_flagp_ms_global=0 sf_flagp_ms_global=0 fs_flagp_ms_global=0 global_mc_flag=1
.param toxn_12_ms_global=0 dxln_12_ms_global=0 dxwn_12_ms_global=0 cjn_12_ms_global=0 cjswn_12_ms_global=0 cjswgn_12_ms_global=0 cgon_12_ms_global=0 cgln_12_ms_global=0 ntoxn_12_ms_global=0 cfn_12_ms_global=0 dvthn_12_ms_global=0 dlvthn_12_ms_global=0 dwvthn_12_ms_global=0 dpvthn_12_ms_global=0 du0n_12_ms_global=0 dlu0n_12_ms_global=0 dwu0n_12_ms_global=0 dpu0n_12_ms_global=0 dvsatn_12_ms_global=0 dlvsatn_12_ms_global=0 dwvsatn_12_ms_global=0 dpvsatn_12_ms_global=0 dk2n_12_ms_global=0 dlk2n_12_ms_global=0 dwk2n_12_ms_global=0 dpk2n_12_ms_global=0 dagsn_12_ms_global=0 dwagsn_12_ms_global=0 dcitn_12_ms_global=0 dlcitn_12_ms_global=0 dwcitn_12_ms_global=0 dpcitn_12_ms_global=0 dpclmn_12_ms_global=0 dlpclmn_12_ms_global=0 dwpclmn_12_ms_global=0 dpua1n_12_ms_global=0 dlucn_12_ms_global=0 dlketan_12_ms_global=0 dwketan_12_ms_global=0 ss_flagn_12_ms_global=0 ff_flagn_12_ms_global=0 monte_flagn_12_ms_global=0 sf_flagn_12_ms_global=0 fs_flagn_12_ms_global=0 toxp_12_ms_global=0 dxlp_12_ms_global=0 dxwp_12_ms_global=0 cjp_12_ms_global=0 cjswp_12_ms_global=0 cjswgp_12_ms_global=0 cgop_12_ms_global=0 cglp_12_ms_global=0 ntoxp_12_ms_global=0 cfp_12_ms_global=0 dvthp_12_ms_global=0 dlvthp_12_ms_global=0 dwvthp_12_ms_global=0 dpvthp_12_ms_global=0 du0p_12_ms_global=0 dlu0p_12_ms_global=0 dwu0p_12_ms_global=0 dpu0p_12_ms_global=0 dvsatp_12_ms_global=0 dwvsatp_12_ms_global=0 dpvsatp_12_ms_global=0 dk2p_12_ms_global=0 dlk2p_12_ms_global=0 dwk2p_12_ms_global=0 dpk2p_12_ms_global=0 dlvoffp_12_ms_global=0 dpvoffp_12_ms_global=0 dagsp_12_ms_global=0 dwagsp_12_ms_global=0 dcitp_12_ms_global=0 dlcitp_12_ms_global=0 dwcitp_12_ms_global=0 dpcitp_12_ms_global=0 deta0p_12_ms_global=0 dpclmp_12_ms_global=0 dua1p_12_ms_global=0 dlucp_12_ms_global=0 dlketap_12_ms_global=0 ss_flagp_12_ms_global=0 ff_flagp_12_ms_global=0 monte_flagp_12_ms_global=0 sf_flagp_12_ms_global=0 fs_flagp_12_ms_global=0 global_mc_flag_12=1
.param toxn_18_ms_global=0 dxln_18_ms_global=0 dxwn_18_ms_global=0 cgon_18_ms_global=0 cgln_18_ms_global=0 cjn_18_ms_global=0 cjswn_18_ms_global=0 cjswgn_18_ms_global=0 cfn_18_ms_global=0 dvthn_18_ms_global=0 dwvthn_18_ms_global=0 dlvthn_18_ms_global=0 dpvthn_18_ms_global=0 du0n_18_ms_global=0 dwu0n_18_ms_global=0 dlu0n_18_ms_global=0 dpu0n_18_ms_global=0 dk2n_18_ms_global=0 dwk2n_18_ms_global=0 dlk2n_18_ms_global=0 dpk2n_18_ms_global=0 dagsn_18_ms_global=0 dwagsn_18_ms_global=0 dvsatn_18_ms_global=0 dwvsatn_18_ms_global=0 dlucn_18_ms_global=0 dlketan_18_ms_global=0 toxp_18_ms_global=0 dxlp_18_ms_global=0 dxwp_18_ms_global=0 cgop_18_ms_global=0 cglp_18_ms_global=0 cjp_18_ms_global=0 cjswp_18_ms_global=0 cjswgp_18_ms_global=0 cfp_18_ms_global=0 dvthp_18_ms_global=0 dwvthp_18_ms_global=0 dlvthp_18_ms_global=0 dpvthp_18_ms_global=0 du0p_18_ms_global=0 dwu0p_18_ms_global=0 dlu0p_18_ms_global=0 dpu0p_18_ms_global=0 dk2p_18_ms_global=0 dwk2p_18_ms_global=0 dlk2p_18_ms_global=0 dpk2p_18_ms_global=0 dagsp_18_ms_global=0 dwagsp_18_ms_global=0 dvsatp_18_ms_global=0 dwvsatp_18_ms_global=0 dlucp_18_ms_global=0 dlketap_18_ms_global=0 ss_flagp_18_ms_global=0 ff_flagp_18_ms_global=0 monte_flagn_18_ms_global=0 monte_flagp_18_ms_global=0 sf_flagp_18_ms_global=0 fs_flagp_18_ms_global=0 global_mc_flag_18=1
.param toxn_18ud15_ms_global=0 dxln_18ud15_ms_global=0 dxwn_18ud15_ms_global=0 cgon_18ud15_ms_global=0 cgln_18ud15_ms_global=0 cjn_18ud15_ms_global=0 cjswn_18ud15_ms_global=0 cjswgn_18ud15_ms_global=0 cfn_18ud15_ms_global=0 dvthn_18ud15_ms_global=0 dwvthn_18ud15_ms_global=0 dlvthn_18ud15_ms_global=0 dpvthn_18ud15_ms_global=0 du0n_18ud15_ms_global=0 dwu0n_18ud15_ms_global=0 dlu0n_18ud15_ms_global=0 dpu0n_18ud15_ms_global=0 dk2n_18ud15_ms_global=0 dwk2n_18ud15_ms_global=0 dlk2n_18ud15_ms_global=0 dpk2n_18ud15_ms_global=0 dagsn_18ud15_ms_global=0 dwagsn_18ud15_ms_global=0 dvsatn_18ud15_ms_global=0 dwvsatn_18ud15_ms_global=0 dlucn_18ud15_ms_global=0 dlketan_18ud15_ms_global=0 toxp_18ud15_ms_global=0 dxlp_18ud15_ms_global=0 dxwp_18ud15_ms_global=0 cgop_18ud15_ms_global=0 cglp_18ud15_ms_global=0 cjp_18ud15_ms_global=0 cjswp_18ud15_ms_global=0 cjswgp_18ud15_ms_global=0 cfp_18ud15_ms_global=0 dvthp_18ud15_ms_global=0 dwvthp_18ud15_ms_global=0 dlvthp_18ud15_ms_global=0 dpvthp_18ud15_ms_global=0 du0p_18ud15_ms_global=0 dwu0p_18ud15_ms_global=0 dlu0p_18ud15_ms_global=0 dpu0p_18ud15_ms_global=0 dk2p_18ud15_ms_global=0 dwk2p_18ud15_ms_global=0 dlk2p_18ud15_ms_global=0 dpk2p_18ud15_ms_global=0 dagsp_18ud15_ms_global=0 dwagsp_18ud15_ms_global=0 dvsatp_18ud15_ms_global=0 dwvsatp_18ud15_ms_global=0 dlucp_18ud15_ms_global=0 dlketap_18ud15_ms_global=0 ss_flagp_18ud15_ms_global=0 ff_flagp_18ud15_ms_global=0 monte_flagn_18ud15_ms_global=0 monte_flagp_18ud15_ms_global=0 sf_flagp_18ud15_ms_global=0 fs_flagp_18ud15_ms_global=0 global_mc_flag_18ud15=1
.param toxn_hvt_ms_global=0 ntoxn_hvt_ms_global=0 dxln_hvt_ms_global=0 dxwn_hvt_ms_global=0 cjn_hvt_ms_global=0 cjswn_hvt_ms_global=0 cjswgn_hvt_ms_global=0 cgon_hvt_ms_global=0 cgln_hvt_ms_global=0 dvthn_hvt_ms_global=0 dlvthn_hvt_ms_global=0 dwvthn_hvt_ms_global=0 dpvthn_hvt_ms_global=0 du0n_hvt_ms_global=0 dlu0n_hvt_ms_global=0 dwu0n_hvt_ms_global=0 dpu0n_hvt_ms_global=0 dvsatn_hvt_ms_global=0 dlvsatn_hvt_ms_global=0 dwvsatn_hvt_ms_global=0 dpvsatn_hvt_ms_global=0 dlvoffn_hvt_ms_global=0 dagsn_hvt_ms_global=0 dwagsn_hvt_ms_global=0 deta0n_hvt_ms_global=0 dpeta0n_hvt_ms_global=0 dk2n_hvt_ms_global=0 dpclmn_hvt_ms_global=0 dua1n_hvt_ms_global=0 dlua1n_hvt_ms_global=0 dpua1n_hvt_ms_global=0 dlatn_hvt_ms_global=0 cfn_hvt_ms_global=0 dpdiblc2n_hvt_ms_global=0 dminvn_hvt_ms_global=0 da0n_hvt_ms_global=0 ss_flagn_hvt_ms_global=0 ff_flagn_hvt_ms_global=0 toxp_hvt_ms_global=0 ntoxp_hvt_ms_global=0 dxlp_hvt_ms_global=0 dxwp_hvt_ms_global=0 cjp_hvt_ms_global=0 cjswp_hvt_ms_global=0 cjswgp_hvt_ms_global=0 cgop_hvt_ms_global=0 cglp_hvt_ms_global=0 dvthp_hvt_ms_global=0 dlvthp_hvt_ms_global=0 dwvthp_hvt_ms_global=0 dpvthp_hvt_ms_global=0 dk2p_hvt_ms_global=0 dleta0p_hvt_ms_global=0 du0p_hvt_ms_global=0 dlu0p_hvt_ms_global=0 dwu0p_hvt_ms_global=0 dpu0p_hvt_ms_global=0 dpclmp_hvt_ms_global=0 dvsatp_hvt_ms_global=0 dlvsatp_hvt_ms_global=0 dwvsatp_hvt_ms_global=0 dpvsatp_hvt_ms_global=0 dagsp_hvt_ms_global=0 dwagsp_hvt_ms_global=0 dpkt1p_hvt_ms_global=0 datp_hvt_ms_global=0 dua1p_hvt_ms_global=0 dlua1p_hvt_ms_global=0 dpua1p_hvt_ms_global=0 cfp_hvt_ms_global=0 dpdiblc2p_hvt_ms_global=0 dminvp_hvt_ms_global=0 dlketap_hvt_ms_global=0 ss_flagp_hvt_ms_global=0 ff_flagp_hvt_ms_global=0 monte_flagn_hvt_ms_global=0 monte_flagp_hvt_ms_global=0 dpvoffn_hvt_ms_global=0 sf_flagn_hvt_ms_global=0 fs_flagn_hvt_ms_global=0 sf_flagp_hvt_ms_global=0 fs_flagp_hvt_ms_global=0 global_mc_flag_hvt=1
.param toxn_lvt_ms_global=0 dxln_lvt_ms_global=0 dxwn_lvt_ms_global=0 cjn_lvt_ms_global=0 cjswn_lvt_ms_global=0 cjswgn_lvt_ms_global=0 cgon_lvt_ms_global=0 cgln_lvt_ms_global=0 ntoxn_lvt_ms_global=0 cfn_lvt_ms_global=0 dvthn_lvt_ms_global=0 dlvthn_lvt_ms_global=0 dwvthn_lvt_ms_global=0 dpvthn_lvt_ms_global=0 du0n_lvt_ms_global=0 dlu0n_lvt_ms_global=0 dwu0n_lvt_ms_global=0 dpu0n_lvt_ms_global=0 dvsatn_lvt_ms_global=0 dlvsatn_lvt_ms_global=0 dwvsatn_lvt_ms_global=0 dpvsatn_lvt_ms_global=0 dk2n_lvt_ms_global=0 dlk2n_lvt_ms_global=0 dwk2n_lvt_ms_global=0 dpk2n_lvt_ms_global=0 dlvoffn_lvt_ms_global=0 dpvoffn_lvt_ms_global=0 dpdiblc2n_lvt_ms_global=0 dagsn_lvt_ms_global=0 dwagsn_lvt_ms_global=0 dleta0n_lvt_ms_global=0 dpclmn_lvt_ms_global=0 dminvn_lvt_ms_global=0 dua1n_lvt_ms_global=0 datn_lvt_ms_global=0 ss_flagn_lvt_ms_global=0 ff_flagn_lvt_ms_global=0 monte_flagn_lvt_ms_global=0 sf_flagn_lvt_ms_global=0 fs_flagn_lvt_ms_global=0 toxp_lvt_ms_global=0 dxlp_lvt_ms_global=0 dxwp_lvt_ms_global=0 cgop_lvt_ms_global=0 cglp_lvt_ms_global=0 cjp_lvt_ms_global=0 cjswp_lvt_ms_global=0 cjswgp_lvt_ms_global=0 cfp_lvt_ms_global=0 dvthp_lvt_ms_global=0 dlvthp_lvt_ms_global=0 dwvthp_lvt_ms_global=0 dpvthp_lvt_ms_global=0 dk2p_lvt_ms_global=0 dlk2p_lvt_ms_global=0 dwk2p_lvt_ms_global=0 dpk2p_lvt_ms_global=0 deta0p_lvt_ms_global=0 dvoffp_lvt_ms_global=0 dlvoffp_lvt_ms_global=0 du0p_lvt_ms_global=0 dlu0p_lvt_ms_global=0 dwu0p_lvt_ms_global=0 dpu0p_lvt_ms_global=0 dpclmp_lvt_ms_global=0 dpdiblc2p_lvt_ms_global=0 dagsp_lvt_ms_global=0 dwagsp_lvt_ms_global=0 ntoxp_lvt_ms_global=0 dvsatp_lvt_ms_global=0 dlvsatp_lvt_ms_global=0 dwvsatp_lvt_ms_global=0 dpvsatp_lvt_ms_global=0 dminvp_lvt_ms_global=0 datp_lvt_ms_global=0 dua1p_lvt_ms_global=0 dlua1p_lvt_ms_global=0 ss_flagp_lvt_ms_global=0 ff_flagp_lvt_ms_global=0 monte_flagp_lvt_ms_global=0 sf_flagp_lvt_ms_global=0 fs_flagp_lvt_ms_global=0 global_mc_flag_lvt=1
.param toxn_na_ms_global=0 dxln_na_ms_global=0 dxwn_na_ms_global=0 cjn_na_ms_global=0 cjswn_na_ms_global=0 cjswgn_na_ms_global=0 cgon_na_ms_global=0 cgln_na_ms_global=0 cfn_na_ms_global=0 dvthn_na_ms_global=0 dlvthn_na_ms_global=0 dwvthn_na_ms_global=0 dpvthn_na_ms_global=0 du0n_na_ms_global=0 dlu0n_na_ms_global=0 dwu0n_na_ms_global=0 dpu0n_na_ms_global=0 dvsatn_na_ms_global=0 dwvsatn_na_ms_global=0 dpdiblc2n_na_ms_global=0 ntoxn_na_ms_global=0 dagsn_na_ms_global=0 dlagsn_na_ms_global=0 dwagsn_na_ms_global=0 dua1n_na_ms_global=0 monte_flagn_na_ms_global=0 ddlcn_na_ms_global=0 global_mc_flag_na=1
.param toxn_na12_ms_global=0 dxln_na12_ms_global=0 dxwn_na12_ms_global=0 cgon_na12_ms_global=0 cgln_na12_ms_global=0 cjn_na12_ms_global=0 cjswn_na12_ms_global=0 cjswgn_na12_ms_global=0 cfn_na12_ms_global=0 dvthn_na12_ms_global=0 dlvthn_na12_ms_global=0 dwvthn_na12_ms_global=0 dpvthn_na12_ms_global=0 du0n_na12_ms_global=0 dlu0n_na12_ms_global=0 dwu0n_na12_ms_global=0 dpu0n_na12_ms_global=0 dvsatn_na12_ms_global=0 dwvsatn_na12_ms_global=0 dk2n_na12_ms_global=0 dlk2n_na12_ms_global=0 dweta0n_na12_ms_global=0 dlcitn_na12_ms_global=0 dpcitn_na12_ms_global=0 datn_na12_ms_global=0 dlatn_na12_ms_global=0 dwatn_na12_ms_global=0 dpatn_na12_ms_global=0 dppdiblc2n_na12_ms_global=0 dlvsatn_na12_ms_global=0 dpvsatn_na12_ms_global=0 ntoxn_na12_ms_global=0 dpclmn_na12_ms_global=0 dwpclmn_na12_ms_global=0 dppclmn_na12_ms_global=0 ff_flagn_na12_ms_global=0 monte_flagn_na12_ms_global=0 ddlcn_na12_ms_global=0 dpdiblc2n_na12_ms_global=0 global_mc_flag_na12=1
.param toxn_na18_ms_global=0 dxln_na18_ms_global=0 dxwn_na18_ms_global=0 cjn_na18_ms_global=0 cjswn_na18_ms_global=0 cjswgn_na18_ms_global=0 cgon_na18_ms_global=0 cgln_na18_ms_global=0 dvthn_na18_ms_global=0 dlvthn_na18_ms_global=0 dwvthn_na18_ms_global=0 dpvthn_na18_ms_global=0 cfn_na18_ms_global=0 du0n_na18_ms_global=0 dlu0n_na18_ms_global=0 dwu0n_na18_ms_global=0 dpu0n_na18_ms_global=0 dvsatn_na18_ms_global=0 dlvsatn_na18_ms_global=0 dwvsatn_na18_ms_global=0 dpvsatn_na18_ms_global=0 dk2n_na18_ms_global=0 dlvoffn_na18_ms_global=0 dppdiblc2n_na18_ms_global=0 dagsn_na18_ms_global=0 dwagsn_na18_ms_global=0 deta0n_na18_ms_global=0 dlk2n_na18_ms_global=0 dwk2n_na18_ms_global=0 dpk2n_na18_ms_global=0 dkt1n_na18_ms_global=0 dlkt2n_na18_ms_global=0 dla0n_na18_ms_global=0 dwa0n_na18_ms_global=0 dlucn_na18_ms_global=0 dlketan_na18_ms_global=0 monte_flagn_na18_ms_global=0 ddlcn_na18_ms_global=0 global_mc_flag_na18=1
.param toxn_na18ud15_ms_global=0 dxln_na18ud15_ms_global=0 dxwn_na18ud15_ms_global=0 cjn_na18ud15_ms_global=0 cjswn_na18ud15_ms_global=0 cjswgn_na18ud15_ms_global=0 cgon_na18ud15_ms_global=0 cgln_na18ud15_ms_global=0 dvthn_na18ud15_ms_global=0 dlvthn_na18ud15_ms_global=0 dwvthn_na18ud15_ms_global=0 dpvthn_na18ud15_ms_global=0 cfn_na18ud15_ms_global=0 du0n_na18ud15_ms_global=0 dlu0n_na18ud15_ms_global=0 dwu0n_na18ud15_ms_global=0 dpu0n_na18ud15_ms_global=0 dvsatn_na18ud15_ms_global=0 dlvsatn_na18ud15_ms_global=0 dwvsatn_na18ud15_ms_global=0 dpvsatn_na18ud15_ms_global=0 dk2n_na18ud15_ms_global=0 dlvoffn_na18ud15_ms_global=0 dppdiblc2n_na18ud15_ms_global=0 dagsn_na18ud15_ms_global=0 dwagsn_na18ud15_ms_global=0 deta0n_na18ud15_ms_global=0 dlk2n_na18ud15_ms_global=0 dwk2n_na18ud15_ms_global=0 dpk2n_na18ud15_ms_global=0 dkt1n_na18ud15_ms_global=0 dlkt2n_na18ud15_ms_global=0 dla0n_na18ud15_ms_global=0 dwa0n_na18ud15_ms_global=0 dlucn_na18ud15_ms_global=0 dlketan_na18ud15_ms_global=0 monte_flagn_na18ud15_ms_global=0 ddlcn_na18ud15_ms_global=0 global_mc_flag_na18ud15=1
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_mac.global nmos ( modelid=1                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag'                 permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=1.95e-009                  toxm=1.95e-009                  dtox=4.06e-010 epsrox=3.9                        wint=0                          lint=0 ll=0                          wl=0                          lln=1 wln=1                          lw=0                          ww=0 lwn=1                          wwn=1                          lwl=0 wwl=0                          llc=0                          wlc=0 lwc=0                          wwc=0                          lwlc=0 wwlc=0                          xl=-4e-009                    xw=6e-009 dlc=5.81e-009                  dwc=0                          xpart=1 toxref=3e-009                     dlcig=2.5e-009                   k1=0.3372 k3=-1                         k3b=0.8                        w0=0 dvt0=0.88                       dvt1=0.79                       dvt2=0.48 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.6                        voffl=0                          dvtp0=1e-006 dvtp1=1.4                        lpe0=0                          lpeb=0 xj=6.7e-008                   ngate=1.476e+020                 ndep=1e+017 nsd=1e+020                     phin=0.13375                    cdsc=0 cdscb=0                          cdscd=0                          nfactor=0.7 ud=0                          lud=0                          wud=0 pud=0                          a1=0                          a2=1 b0=0                          b1=0                          dwg=0 dwb=0                          pdiblc1=0                          pdiblcb=1 drout=0.56                       pvag=2                          delta=0.01 pscbe1=1e+009                     pscbe2=1e-020                     fprout=78 pdits=0.0027                     pditsd=0                          pditsl=0 rsh=18.0                       rdsw=120                        rsw=0 rdw=0                          prwg=0                          prwb=0 wr=1                          alpha0=1e-008                     alpha1=1.5 beta0=12                         agidl=1e-006                     bgidl=3.459e+009 cgidl=0.295                      egidl=0.27814                    bigbacc=0.0074708 cigbacc=0.2809                     nigbacc=4.05                       aigbinv=0.2415 bigbinv=0.0309                     cigbinv=0.006                      eigbinv=1.1 nigbinv=1                          bigc=0.00159                    cigc=1e-005 cigsd=2e-020                     nigc=3.083                      poxedge=1 pigcd=2.46                       ntox=1                          xrcrg1=12 xrcrg2=1                          vfbsdoff=0.01                       lvfbsdoff=0 wvfbsdoff=0                          pvfbsdoff=0                          cgso=8.14e-011 cgdo=8.14e-011                  cgbo=0                          cgdl=2.4209e-011 cgsl=2.4209e-011                clc=0                          cle=0.6 cf='6.62e-011+9.73e-11*ccoflag'                                       ckappas=0.6 ckappad=0.6                        acde=0.3                        moin=6.5 noff=2.5                        voffcv=-0.098559                  tvfbsdoff=0.1 ltvfbsdoff=0                          wtvfbsdoff=0                          ptvfbsdoff=0 kt1l=0                          ute=-1                         prt=0 fnoimod=1.000000e+00               tnoimod=1                          em=1.000000e+06 ef=9.000000e-01               noia=0                          noib=0 noic=0                          lintnoi=-2.790000e-08              jss=4.32e-07 jsd=4.32e-07                   jsws=1.17e-13                   jswd=1.17e-13 jswgs=1.17e-13                   jswgd=1.17e-13                   njs=1.03 njd=1.03                       ijthsfwd=0.01                       ijthdfwd=0.01 ijthsrev=0.01                       ijthdrev=0.01                       bvs=8.219999 bvd=8.219999                   xjbvs=1                          xjbvd=1 njtsswg=16                         xtsswgs=0.16                       xtsswgd=0.16 tnjtsswg=1                          vtsswgs=1                          vtsswgd=1 pbs=0.672                      pbd=0.672                      cjs=0.001428 cjd=0.001428                   mjs=0.321                      mjd=0.321 pbsws=0.480                      pbswd=0.480                      cjsws=1.069e-010 cjswd=1.069e-010                 mjsws=0.016                      mjswd=0.016 pbswgs=0.990                      pbswgd=0.990                      cjswgs=2.9e-010 cjswgd=2.9e-010                   mjswgs=0.725                      mjswgd=0.725 tpb=0.00114                    tcj=0.00072                    tpbsw=0.00244 tcjsw=0.00020                    tpbswg=0.00171                    tcjswg=0.00124 xtis=3                          xtid=3                          dmcg=3.8e-008 dmci=3.8e-008                   dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=2.64e-009 rshg=16.42                      gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          lnfactor=0 pnfactor=0                          wnfactor=0                          pk2we=0 lk2we=0                          wk2we=0                          k2we=0.0000 pku0we=-1e-18                     wku0we=3e-11                      lku0we=4.5e-11 ku0we=-0.0016                    pkvth0we=1.3e-018                   wkvth0we=-4.1e-011 lkvth0we=-1.05e-011                 kvth0we=0.00053                    wec=-9093.6 web=2153.1                     scref=1e-6                       rnoia=0 rnoib=0                          tnoia=0                          wpemod=1 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.2                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.4 bidirectionflag='bidirectionflag_mos' iboffn_flag='iboffn_flag' iboffp_flag='iboffp_flag' sigma_factor='sigma_factor' ccoflag='ccoflag' rcoflag='rcoflag' rgflag='rgflag' mismatchflag='mismatchflag_mos' globalflag='globalflag_mos' totalflag='totalflag_mos' designflag='designflag_mos' global_factor='global_factor' local_factor='local_factor' sigma_factor_flicker='sigma_factor_flicker' noiseflag='noiseflagn' noiseflag_mc='noiseflagn_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w1='2.3875*0.35355' w2='0.70711*-0.35355' w3='0.54772*-0.0052117' w4='0.54772*-0.40307' w5='0.54772*-0.64548' w6='0.54772*-0.049915' w7='0.54772*-0.11513' w8='0.54772*-0.39385' w9='0' w10='0' tox_c='toxn'                     dxl_c='dxln'                     dxw_c='dxwn' cj_c='cjn'                      cjsw_c='cjswn'                    cjswg_c='cjswgn' cgo_c='cgon'                     cgl_c='cgln'                     ddlc_c='ddlcn' cf_c='cfn'                      ntox_c='ntoxn'                    dvth_c='dvthn' dlvth_c='dlvthn'                   dwvth_c='dwvthn'                   dpvth_c='dpvthn' du0_c='du0n'                     dlu0_c='dlu0n'                    dwu0_c='dwu0n' dpu0_c='dpu0n'                    dvsat_c='dvsatn'                   dlvsat_c='dlvsatn' dwvsat_c='dwvsatn'                  dpvsat_c='dpvsatn'                  dk2_c='dk2n' dlk2_c='dlk2n'                    dwk2_c='dwk2n'                    dpk2_c='dpk2n' dvoff_c='dvoffn'                   dlvoff_c='dlvoffn'                  dwvoff_c='dwvoffn' dpvoff_c='dpvoffn'                  dpdiblc2_c='dpdiblc2n'                dlpdiblc2_c='dlpdiblc2n' dwpdiblc2_c='dwpdiblc2n'               dppdiblc2_c='dppdiblc2n'               dags_c='dagsn' dlags_c='dlagsn'                   dwags_c='dwagsn'                   dpags_c='dpagsn' dnfactor_c='dnfactorn'                dlnfactor_c='dlnfactorn'               dwnfactor_c='dwnfactorn' dpnfactor_c='dpnfactorn'               dcit_c='dcitn'                    dlcit_c='dlcitn' dwcit_c='dwcitn'                   dpcit_c='dpcitn'                   deta0_c='deta0n' dleta0_c='dleta0n'                  dweta0_c='dweta0n'                  dpeta0_c='dpeta0n' dpclm_c='dpclmn'                   dlpclm_c='dlpclmn'                  dwpclm_c='dwpclmn' dppclm_c='dppclmn'                  jtsswg_c='jtsswgn'                  dminv_c='dminvn' dketa_c='dketan'                   dlketa_c='dlketan'                  dwketa_c='dwketan' dpketa_c='dpketan'                  dua1_c='dua1n'                    dlua1_c='dlua1n' dwua1_c='dwua1n'                   dpua1_c='dpua1n'                   dat_c='datn' dlat_c='dlatn'                    dwat_c='dwatn'                    dpat_c='dpatn' ss_flag_c='ss_flagn'                 ff_flag_c='ff_flagn'                 sf_flag_c='sf_flagn' fs_flag_c='fs_flagn'                 monte_flag_c='monte_flagn'             c1f_c='c1fn' c2f_c='c2fn'                     c3f_c='c3fn' global_mc='global_mc_flag' tox_g='toxn_ms_global'           dxl_g='dxln_ms_global'           dxw_g='dxwn_ms_global' cj_g='cjn_ms_global'            cjsw_g='cjswn_ms_global'          cjswg_g='cjswgn_ms_global' cgo_g='cgon_ms_global'           cgl_g='cgln_ms_global'           cf_g='cfn_ms_global' ntox_g='ntoxn_ms_global'          dvth_g='dvthn_ms_global'          dlvth_g='dlvthn_ms_global' dwvth_g='dwvthn_ms_global'         dpvth_g='dpvthn_ms_global'         du0_g='du0n_ms_global' dlu0_g='dlu0n_ms_global'          dwu0_g='dwu0n_ms_global'          dpu0_g='dpu0n_ms_global' dvsat_g='dvsatn_ms_global'         dlvsat_g='dlvsatn_ms_global'        dwvsat_g='dwvsatn_ms_global' dpvsat_g='dpvsatn_ms_global'        dk2_g='dk2n_ms_global'           dlk2_g='dlk2n_ms_global' dwk2_g='dwk2n_ms_global'          dlvoff_g='dlvoffn_ms_global'        dpvoff_g='dpvoffn_ms_global' dpdiblc2_g='dpdiblc2n_ms_global'      dppdiblc2_g='dppdiblc2n_ms_global'     dags_g='dagsn_ms_global' dwags_g='dwagsn_ms_global'         dlcit_g='dlcitn_ms_global'         dpcit_g='dpcitn_ms_global' dpclm_g='dpclmn_ms_global'         dminv_g='dminvn_ms_global'         dketa_g='dketan_ms_global' dlketa_g='dlketan_ms_global'        dpketa_g='dpketan_ms_global'        dua1_g='dua1n_ms_global' dat_g='datn_ms_global'           ss_flag_g='ss_flagn_ms_global'       ff_flag_g='ff_flagn_ms_global' monte_flag_g='monte_flagn_ms_global'   deta0_g='deta0n_ms_global'         sf_flag_g='sf_flagn_ms_global' fs_flag_g='fs_flagn_ms_global' weight1=-3.2637736 weight2=1.9622013 weight3=-1.3576101 weight4=-0.62893082 weight5=-0.43842138 tox_1=4.0248948e-012 tox_2=-9.9546871e-012 tox_3=1.2167984e-013 tox_4=3.7476951e-011 tox_5=7.2868905e-013 dxl_1=9.1129882e-011 dxl_2=-2.2538971e-010 dxl_3=2.7548964e-012 dxl_4=-8.485289e-010 dxl_5=1.6498979e-011 dxw_1=-6.912291e-010 dxw_2=-7.9677896e-010 dxw_3=-5.351993e-011 dxw_4=-5.6696926e-025 dxw_5=-5.9028923e-009 cj_1=9.4466e-006 cj_2=-3.0912e-006 cj_3=5.1272e-007 cj_4=-1.3389e-021 cj_5=-7.3543e-007 cjsw_1=7.0717e-013 cjsw_2=-2.3141e-013 cjsw_3=3.8382e-014 cjsw_4=-1.4248e-029 cjsw_5=-5.5054e-014 cjswg_1=1.9184e-012 cjswg_2=-6.2777e-013 cjswg_3=1.0412e-013 cjswg_4=4.0403e-028 cjswg_5=-1.4935e-013 cgo_1=-5.3848e-013 cgo_2=1.7621e-013 cgo_3=-2.9227e-014 cgo_4=9.673e-029 cgo_5=4.1921e-014 cgl_1=-1.6015e-013 cgl_2=5.2406e-014 cgl_3=-8.6922e-015 cgl_4=3.2268e-030 cgl_5=1.2468e-014 cf_1=-4.3793e-013 cf_2=1.433e-013 cf_3=-2.3769e-014 cf_4=8.8236e-030 cf_5=3.4093e-014 ntox_1=-0.018901 ntox_2=0.0061849 ntox_3=-0.0010259 ntox_4=1.6805e-017 ntox_5=0.0014714 dvth_1=0.0031311 dvth_2=0.0040311 dvth_3=-0.00018211 dvth_4=1.7396e-018 dvth_5=-0.00084981 dlvth_1=6.6819e-011 dlvth_2=9.043e-011 dlvth_3=1.4159e-011 dlvth_4=-2.2585e-026 dlvth_5=-1.8507e-011 dwvth_1=2.3252e-010 dwvth_2=5.3451e-011 dwvth_3=-2.0771e-011 dwvth_4=3.0823e-025 dwvth_5=-3.0027e-011 dpvth_1=2.1586e-017 dpvth_2=1.6912e-017 dpvth_3=1.9847e-018 dpvth_4=3.1216e-033 dpvth_5=-4.3306e-018 du0_1=0.00012295 du0_2=0.00024165 du0_3=3.6177e-005 du0_4=-7.2484e-020 du0_5=-4.7951e-005 dlu0_1=-6.1084e-013 dlu0_2=5.6833e-012 dlu0_3=4.3492e-013 dlu0_4=-2.7602e-027 dlu0_5=-7.333e-013 dwu0_1=8.1582e-012 dwu0_2=1.3962e-011 dwu0_3=-2.1138e-012 dwu0_4=-4.5445e-027 dwu0_5=-2.5495e-012 dpu0_1=4.4097e-019 dpu0_2=5.3538e-018 dpu0_3=-2.5756e-019 dpu0_4=3.8918e-034 dpu0_5=-1.1893e-018 dvsat_1=1158.2 dvsat_2=-378.55 dvsat_3=11.779 dvsat_4=1.2538e-012 dvsat_5=-89.735 dlvsat_1=6.9637e-006 dlvsat_2=5.8878e-005 dlvsat_3=7.6832e-007 dlvsat_4=4.1677e-020 dlvsat_5=-8.0822e-006 dwvsat_1=2.4601e-005 dwvsat_2=-7.621e-006 dwvsat_3=-4.8725e-005 dwvsat_4=7.1567e-021 dwvsat_5=-1.4928e-006 dpvsat_1=3.6065e-012 dpvsat_2=3.067e-011 dpvsat_3=-2.8384e-012 dpvsat_4=-6.2663e-027 dpvsat_5=-5.9883e-012 dk2_1=0.00087071 dk2_2=0.0011775 dk2_3=0.00057452 dk2_4=-1.7426e-019 dk2_5=-0.00024905 dlk2_1=9.2454e-012 dlk2_2=-3.2005e-012 dlk2_3=2.0935e-011 dlk2_4=1.6293e-026 dlk2_5=-8.9218e-013 dwk2_1=1.8491e-011 dwk2_2=-6.401e-012 dwk2_3=4.1869e-011 dwk2_4=5.1577e-027 dwk2_5=-1.7844e-012 dlvoff_1=-7.4926e-012 dlvoff_2=2.3159e-012 dlvoff_3=1.5449e-011 dlvoff_4=7.5669e-027 dlvoff_5=4.4951e-013 dpvoff_1=1.3035e-018 dpvoff_2=-4.0289e-019 dpvoff_3=-2.6877e-018 dpvoff_4=-1.4638e-033 dpvoff_5=-7.8201e-020 dpdiblc2_1=-2.8351e-005 dpdiblc2_2=9.2773e-006 dpdiblc2_3=-1.5388e-006 dpdiblc2_4=1.5825e-020 dpdiblc2_5=2.2072e-006 dppdiblc2_1=-7.5603e-019 dppdiblc2_2=2.474e-019 dppdiblc2_3=-4.1034e-020 dppdiblc2_4=-2.6217e-034 dppdiblc2_5=5.8858e-020 dags_1=0.050169 dags_2=0.045072 dags_3=-0.017476 dags_4=3.2926e-017 dags_5=-0.011951 dwags_1=1.0367e-009 dwags_2=3.0556e-009 dwags_3=-3.2371e-010 dwags_4=3.8482e-025 dwags_5=-3.5432e-010 dlcit_1=2.8761e-013 dlcit_2=-9.0612e-014 dlcit_3=-3.9305e-013 dlcit_4=7.5835e-029 dlcit_5=-1.8943e-014 dpcit_1=-1.6795e-019 dpcit_2=5.2767e-020 dpcit_3=2.463e-019 dpcit_4=-1.6862e-034 dpcit_5=1.0919e-020 dpclm_1=-0.011813 dpclm_2=0.0038656 dpclm_3=-0.00064116 dpclm_4=2.0595e-017 dpclm_5=0.00091965 dminv_1=-0.0070878 dminv_2=0.0023193 dminv_3=-0.0003847 dminv_4=1.2357e-017 dminv_5=0.00055179 dketa_1=-0.0018901 dketa_2=0.00061849 dketa_3=-0.00010259 dketa_4=3.7416e-018 dketa_5=0.00014714 dlketa_1=-2.0217e-010 dlketa_2=7.106e-011 dlketa_3=-5.8309e-010 dlketa_4=-3.027e-025 dlketa_5=2.0567e-011 dpketa_1=-2.7736e-017 dpketa_2=9.6015e-018 dpketa_3=-6.2804e-017 dpketa_4=-2.9117e-033 dpketa_5=2.6765e-018 dua1_1=1.8901e-012 dua1_2=-6.1849e-013 dua1_3=1.0259e-013 dua1_4=3.1296e-028 dua1_5=-1.4714e-013 dat_1=1606.6 dat_2=-525.72 dat_3=87.198 dat_4=1.1874e-012 dat_5=-125.07 ss_flag_1=0.046227 ss_flag_2=-0.016003 ss_flag_3=0.10467 ss_flag_4=-1.4034e-018 ss_flag_5=-0.0044609 ff_flag_1=-0.048277 ff_flag_2=0.014922 ff_flag_3=0.099544 ff_flag_4=-8.7429e-017 ff_flag_5=0.0028963 monte_flag_1=0.0759417 monte_flag_2=-0.187825 monte_flag_3=0.00229575 monte_flag_4=-0.707108 monte_flag_5=0.0137492 sigma_local=1                          a_1=0.95976 b_1=-0.00265699                c_1=-0.00151863                d_1=0.000362349 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1.04934                    b_2=-0.00148031                c_2=-0.00335035 d_2=-0.000662885               a_3=1.00581                    b_3=-0.00534195 c_3=-0.00573488                d_3=-0.000284785               e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.84 b_4=-0.00095                   c_4=-0.004                     d_4=0.00002 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=0.82                       b_5=-0.00475                   c_5=0.001 d_5=-0.00018                   e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.004                      mis_a_2=0.15                       mis_a_3=0.15 mis_b_1=0.003                      mis_b_2=0.1                        mis_b_3=0 mis_c_1=0.7                        mis_c_2=0                          mis_c_3=0 mis_d_1=0.00085                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.005                      mis_e_2=0.06                       mis_e_3=0.08 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-4e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0 cf0=6.62e-011                  cco=9.73e-11 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.49                       l_rjtsswg=2.5e-5                     ll_rjtsswg=3 w_rjtsswg=0                          ww_rjtsswg=0                          p_rjtsswg=0 noimod=6                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718                      tnoiamax=8273641.5175 tnoiac1=1759434.0988               tnoiac2=128113.2824                rnoiamax=0.4186 rnoiac1=0.0097201                  rnoiac2=0.3736 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6                sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=0                   lreflod=1e-6                llodref=3 lod_clamp=-1e90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=1 kvth00=0                   lkvth00=0                   wkvth00=0 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=0                   lku000=0                   wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0                   lkvth000=0                   wkvth000=0         		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=0                   wku01=0 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=0                   wkvth01=0 pkvth01=0                   llodvth1=1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.06               lku02=1.5e-7              wku02=7e-8 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=-0.5 kvth02=7e-3                lkvth02=-9e-9               wkvth02=16e-9 pkvth02=1e-15               llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=-0.03               lku03=7e5                 wku03=-5e-8 pku03=0                   tku03=0                   llodku03=-1 wlodku03=1                   kvsat3=0 kvth03=9e-3                lkvth03=-3e-9               wkvth03=-2e-8 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=-0.000                   lku003=-0.0e-9                   wku003=-0e-9         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0.0e-3                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='0.15*01'           wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl='1.4e-12*1'         ldplkvth0=1.5                 pkvth0dpl=0.0e-19 ku0dpl='0.50*1'            wku0dpl=7e-8                wdplku0=1 lku0dpl=11.0e-8              ldplku0=1.0                 pku0dpl=0.0e-11 keta0dpl='0.07*0'            wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0.00                wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx='0.25*1'            wku0dpx=0e-9                wdpxku0=1 lku0dpx='1.0e-8*1'          ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps='0.1*1'             wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='-0.70*1'           wku0dps=-0.0e-9             wdpsku0=1 lku0dps='9.0e-15*1'         ldpsku0=2.0                 pku0dps='-7.0e-23*0' keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps='-0.3*0'            wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa='0.01*0'            wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa='1.0e-9*0'          ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa='0.050*0'           wku0dpa=0e-7                wdpaku0=1 lku0dpa=0.0e-11             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=-0.0                wka0dpa=0                   wdpaka0=1 lka0dpa=-0.0e-7             ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa='1.5*0'             wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2='0.005*1'           wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2='3e-9*1'            ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.000               wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2='2.5e-5*1'          ldp2ku0=0.5                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2='0.5*0'             wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx='0.050*2'           wkvth0enx='8.0e-9*1'          wenxkvth0=1 lkvth0enx='1.0e-8*1'          lenxkvth0=1.0                 pkvth0enx=0 ku0enx='-0.90*1.7'         wku0enx='-0.9e-8*1.5'       wenxku0=1 lku0enx='2.0e-7*1'          lenxku0=1.0                 pku0enx='-3.0e-16*1.7' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0.0                 wka0enx=0                   wenxka0=1 lka0enx='1.0e-7*2'          lenxka0=1.0                 pka0enx='1.0e-14*1.7' kvsatenx=-0.0                wenx=0                   ku0enx0='0.15*0' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.01e-6 kvth0eny='0.04*1.7'          wkvth0eny='4.0e-10*4'         wenykvth0=1 lkvth0eny='1.0e-7*1.7'        lenykvth0=1.0                 pkvth0eny=0 ku0eny='-0.70*2'           wku0eny='-1.1e-8*1'         wenyku0=1 ku0eny0='0.025*0'           wku0eny0=0                   weny0ku0=1 lku0eny='6.0e-10*1.7'       lenyku0=1.5                 pku0eny=-0.0e-14 keta0eny=0.00                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-8             wenyka0=1 lka0eny='-6.0e-8*1.7'       lenyka0=1.0                 pka0eny='1.0e-14*1.7' kvsateny=-0.0                weny=0 kvth0eny1=0.000              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=0 ku0eny1='0.15*1.7'         wku0eny1=0.0e-8             weny1ku0=1 lku0eny1='1.0e-5*1.0'       leny1ku0=1.0                pku0eny1=-0.0e-14 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1.0                pka0eny1=0 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=-0.045              wkvth0rx=-0.0e-5             wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0.0e-16 ku0rx='0.3'               wku0rx=0.0e-8              wrxku0=1.0 lku0rx='-3.5e-10*0'        lrxku0=1                   pku0rx=0.0e-15 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.0                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=0.9027e-5           ringymin=0.117e-6 kvth0ry='-0.03*1'           wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry=0.0e-8              lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry='-0.02*1'           wku0ry=-0.0e-8             wryku0=1.0 lku0ry='-1.0e-8*1'         lryku0=1.0                 pku0ry=-0.0e-16 keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry=0                   wry=0 kvth0ry0=0.01                ku0ry0=0.02 sfxref=9.0e-8            sfxmax=3.906e-6           minwodx=0.0e-6 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0009            lkvth0odx1b=0.0e-7            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.0028           lku0odx1b=0.8e-10           lodx1bku0=1.0 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6              sfymax=10e-6             minwody=0.9e-6 wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-1.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.000            lkvth0odyb=0.0e-10           lodybkvth0=1.0 wkvth0odyb=-2.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.03             lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-1.0e-7           wodybku0=1.0               pku0odyb=0 web_mac=0  wec_mac=0 kvsatwe=0.0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_mac.1 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=9.01e-06                   vth0=0.3801863 lvth0=1.6766525e-009             wvth0=-2.69231e-008              pvth0=-1.5178598e-015 k2=-0.014561973               lk2=-9.4171827e-014            wk2=-6.5204909e-009 pk2=-5.8841761e-020            minv=-0.42453                   cit=0.0011899043 wcit=-1.7205329e-010            voff=-0.1566818                 lvoff=-2.409094e-008 wvoff=5.186393e-009              pvoff=-3.2832359e-015            eta0=0.0096711111 weta0=-6.0440267e-009            etab=-0.034548457               wetab=-9.5406724e-009 u0=0.018409273                wu0=3.8480303e-010             ua=-1.6009732e-009 lua=4.282724e-017              wua=1.032247e-016              pua=-6.6227134e-023 ub=1.983289e-018              wub=-9.0861868e-026            uc=1.8646376e-010 luc=-3.802364e-017             wuc=-1.8363892e-017            puc=-1.603864e-023 vsat=132796.3                   wvsat=-0.025183444               a0=2.2936034 la0=-4.4256733e-007            wa0=5.7953013e-009             pa0=4.00966e-013 ags=1.1901392                  lags=1.0688401e-006             wags=-7.7878351e-008 pags=8.8741184e-014             keta=-0.014753628               lketa=-7.7382942e-008 wketa=3.2448713e-008             pketa=-2.00483e-014              pclm=0.4 lpclm=1.1130524e-015             wpclm=1.1142896e-015             ppclm=-1.002415e-020 pdiblc2=0.00051237275              lpdiblc2=-1.1130524e-010            wpdiblc2=-1.1142897e-010 ppdiblc2=1.002415e-015              aigbacc=0.013223093                waigbacc=-1.2692456e-010 aigc=0.010827522                laigc=-3.3772635e-011            waigc=7.5769128e-011 paigc=-9.0077012e-019            aigsd=0.0096880559               laigsd=6.6932764e-011 waigsd=2.2098242e-011             paigsd=3.6594062e-018             bigsd=0.00050424727 wbigsd=-3.8480303e-012            tvoff=0.00251219                 ltvoff=-3.46739e-010 wtvoff=-1.6168e-010               ptvoff=1.06044e-016               kt1=-0.1617 lkt1=-1.0172267e-014            wkt1=4.6800167e-013             pkt1=-4.210143e-018 kt2=-0.070615243               wkt2=1.015195e-008              ua1=1.5947215e-009 lua1=-4.1553233e-017            wua1=-5.5076454e-017            pua1=3.6439189e-024 ub1=-1.3716307e-018            wub1=4.1703784e-026             uc1=1.0961448e-010 luc1=-3.450433e-017             wuc1=-2.6814585e-018            puc1=9.6231841e-024 at=130000                     jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=0 pcit=0                          lu0=0                          pu0=0 lat=0                          lvsat=0                          pvsat=0 wat=0                          pat=0                          leta0=0 peta0=0                          vth0_mcl=9.93715e-05                lvth0_mcl=1.11155e-10 wvth0_mcl=-8.95934e-10               pvth0_mcl=-1.00217e-15               u0_mcl=3.72169e-06 wu0_mcl=-3.35547e-11               a0_sf=0.0116652                  la0_sf=-1.05057e-07 wa0_sf=-5.56391e-09               pa0_sf=5.01086e-14                lu0_mcl=-3.33463e-12 pu0_mcl=3.0065e-17 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.2 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.38799684 lvth0=-5.3215902e-009            wvth0=-3.1831443e-008            pvth0=2.8800157e-015 k2=-0.015581493               lk2=9.1339634e-010             wk2=-2.6189797e-009 pk2=-3.4958128e-015            minv=-0.42453                   cit=0.00043135249 wcit=-7.4193069e-010            voff=-0.1779059                 lvoff=-5.074142e-009 wvoff=-2.6196974e-009            pvoff=3.7110211e-015             eta0=0.0096711111 weta0=-6.0440267e-009            etab=-0.034548457               wetab=-9.5406724e-009 u0=0.018352271                wu0=3.2689678e-010             ua=-1.4761759e-009 lua=-6.8991176e-017            wua=5.942712e-017              pua=-2.6984503e-023 ub=2.0089136e-018             wub=-1.3419172e-025            uc=1.4313981e-010 luc=7.9462737e-019             wuc=-2.8277091e-017            puc=-7.1564141e-024 vsat=132796.3                   wvsat=-0.025183444               a0=1.556771 la0=2.1763449e-007             wa0=1.3019281e-006             pa0=-7.60369e-013 ags=1.6196044                  lags=6.8403929e-007             wags=5.1811237e-007 pags=-4.452665e-013             keta=-0.081615889               lketa=-1.7474356e-008 wketa=-3.4534404e-008            pketa=3.9968573e-014             pclm=0.25385025 lpclm=1.3095018e-007             wpclm=-9.2075009e-008            ppclm=8.2499199e-014 pdiblc2=-0.00015175045             lpdiblc2=4.8374915e-010             wpdiblc2=1.4066912e-009 ppdiblc2=-3.578207e-016             aigbacc=0.013091601                waigbacc=-1.2093426e-010 aigc=0.010786213                laigc=3.2400783e-012             waigc=8.8573946e-011 paigc=-1.2373887e-017            aigsd=0.0097959832               laigsd=-2.9770148e-011 waigsd=5.1627786e-011             paigsd=-2.2799065e-017            bigsd=0.00050308688 wbigsd=6.6024758e-012             tvoff=0.00208874                 ltvoff=3.26697e-011 wtvoff=9.57373e-011               ptvoff=-1.24601e-016              kt1=-0.16179387 lkt1=8.4096204e-011             wkt1=1.0744208e-008             pkt1=-9.6306011e-015 kt2=-0.071512774               wkt2=1.1683471e-008             ua1=1.945523e-009 lua1=-3.5587134e-016            wua1=-1.0323302e-016            pua1=4.6792205e-023 ub1=-1.6527444e-018            wub1=1.18779e-025               uc1=5.2586825e-011 luc1=1.6592451e-017             wuc1=3.201991e-017              puc1=-2.1469242e-023 at=139911.11                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=6.7966242e-010 pcit=5.1061015e-016             lu0=5.1073227e-011             pu0=5.1884002e-017 lub=-2.29596e-026              pub=3.8823547e-032             laigbacc=1.1781666e-010 paigbacc=-5.3673106e-018            lbigsd=1.0397128e-012             pbigsd=-9.3636535e-018 lkt2=8.041879e-010              pkt2=-1.3722424e-015            lub1=2.5187793e-025 pub1=-6.9059396e-032            lat=-0.0088803556              lvsat=0 pvsat=0                          wat=0                          pat=0 leta0=0                          peta0=0                          vth0_mcl=0.00044487 lvth0_mcl=-1.98412e-10               wvth0_mcl=-4.01095e-09               pvth0_mcl=1.78888e-15 a0_sf=-0.210233                  la0_sf=9.37639e-08                wa0_sf=1.00273e-07 pa0_sf=-4.47221e-14               ags_ss=-0.0792889                 ags_ff=0.118933 ags_sf=-0.0495556                 ags_fs=0.0594666                  lags_ss=7.10428e-08 lags_ff=-1.06564e-07               lags_sf=4.44018e-08                lags_fs=-5.32821e-08 wags_ss=1.4e-14                    wags_ff=1.8e-13                    wags_sf=9e-15 wags_fs=-1.1e-14                   pags_ss=-3.6e-20                   pags_ff=1e-19 pags_sf=4e-20                      pags_fs=-4.8e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.3 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.38929891 lvth0=-5.9023129e-009            wvth0=-3.3582934e-008            pvth0=3.6611806e-015 k2=-0.015662817               lk2=9.4966664e-010             wk2=-7.2072926e-009 pk2=-1.4494253e-015            minv=-0.42453                   cit=0.0015254332 wcit=1.9430771e-010             voff=-0.18828204                lvoff=-4.4638158e-010 wvoff=1.3087748e-008             pvoff=-3.2944994e-015            eta0=0.0096711111 weta0=-6.0440267e-009            etab=-0.034548457               wetab=-9.5406724e-009 u0=0.018400167                wu0=2.7621718e-010             ua=-1.5650944e-009 lua=-2.9333506e-017            wua=8.0679368e-018             pua=-4.0783072e-024 ub=2.0684664e-018             wub=-4.513562e-026             uc=1.7230364e-010 luc=-1.2212443e-017            wuc=-4.6148124e-017            puc=8.1406668e-025 vsat=147906.08                  wvsat=-0.038872907               a0=2.9153365 la0=-3.8828569e-007            wa0=-5.3503842e-007            pa0=5.8918076e-014 ags=3.3726991                  lags=-9.7840955e-008            wags=-8.240719e-007 pags=1.5334768e-013             keta=-0.10844576                lketa=-5.5082326e-009 wketa=6.8854654e-008             pketa=-6.1429472e-015            pclm=0.15471424 lpclm=1.7516484e-007             wpclm=2.1902235e-008             ppclm=3.1665348e-014 pdiblc2=0.00096328965              lpdiblc2=-1.3558739e-011            wpdiblc2=3.3061342e-010 ppdiblc2=1.2211e-016                aigbacc=0.013501499                waigbacc=-3.6842734e-010 aigc=0.010779911                laigc=6.0510222e-012             waigc=8.4702583e-011 paigc=-1.064726e-017             aigsd=0.0097471722               laigsd=-8.0004219e-012 waigsd=-4.88406e-011              paigsd=2.2009835e-017             bigsd=0.00056139071 wbigsd=-6.6294403e-011            tvoff=0.00220832                 ltvoff=-2.06619e-011 wtvoff=-3.45722e-011              ptvoff=-6.64832e-017              kt1=-0.14789643 lkt1=-6.1141608e-009            wkt1=-9.275929e-009             pkt1=-7.0162006e-016 kt2=-0.074238567               wkt2=1.2709882e-008             ua1=1.4683811e-009 lua1=-1.4306603e-016            wua1=-1.3247317e-016            pua1=5.983331e-023 ub1=-1.3025272e-018            wub1=3.7568361e-026             uc1=1.3733024e-010 luc1=-2.1203114e-017            wuc1=-5.2622637e-017            puc1=1.6281334e-023 at=154489.99                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.9170243e-010 pcit=9.3047822e-017             lu0=2.9711597e-011             pu0=7.4487101e-017 lub=-4.9520166e-026            pub=-8.9547335e-034            laigbacc=-6.4997541e-011 paigbacc=1.050146e-016              lbigsd=-2.4963795e-011            pbigsd=2.3148354e-017 lkt2=2.0198917e-009             pkt2=-1.8300219e-015            lub1=9.5681051e-026 pub1=-3.283945e-032             lat=-0.015382536               lvsat=-0.0067389626 pvsat=6.1055001e-009             wat=0.014303006                pat=-6.3791407e-009 leta0=0                          peta0=0                          ags_ss=0.0981197 ags_ff=-0.156239                  ags_sf=0.0681193                  ags_fs=-0.0781191 lags_ss=-8.08138e-09               lags_ff=1.61627e-08                lags_sf=-8.08135e-09 lags_fs=8.08136e-09                wags_ss=4.44e-13                   wags_ff=7.08e-13 wags_sf=-2.8e-14                   wags_fs=2.04e-13                   pags_ss=-2.9e-20 pags_ff=-2.8e-20                   pags_sf=-1.4e-20                   pags_fs=-1.4e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.4 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.36985536 lvth0=-1.7802816e-009            wvth0=-1.8276777e-008            pvth0=4.1627547e-016 k2=-0.012210364               lk2=2.177466e-010              wk2=-1.137847e-008 pk2=-5.6513573e-016            minv=-0.42453                   cit=0.0013809444 wcit=1.0053135e-009             voff=-0.18176071                lvoff=-1.8289053e-009 wvoff=1.8545258e-009             pvoff=-9.1305633e-016            eta0=0.0096711111 weta0=-6.0440267e-009            etab=-0.034548421               wetab=-9.5409825e-009 u0=0.018777472                wu0=6.1244538e-010             ua=-1.7720854e-009 lua=1.4548594e-017             wua=-3.7312989e-017            pua=5.5424491e-024 ub=2.011493e-018              wub=-2.0207516e-026            uc=1.2833947e-010 luc=-2.8920389e-018            wuc=-2.9932323e-017            puc=-2.6236832e-024 vsat=115442.74                  wvsat=-0.016072248               a0=3.1721562 la0=-4.4273148e-007            wa0=-1.575924e-008             pa0=-5.116911e-014 ags=2.9240719                  lags=-2.7319918e-009            wags=-2.1679188e-007 pags=2.4604318e-014             keta=-0.06385227                lketa=-1.4962053e-008 wketa=1.8968778e-008             pketa=4.4328585e-015             pclm=0.90429693 lpclm=1.6253308e-008             wpclm=2.4691079e-007             ppclm=-1.6036465e-014 pdiblc2=0.00092234931              lpdiblc2=-4.8793863e-012            wpdiblc2=7.0023724e-010 ppdiblc2=4.3749753e-017             aigbacc=0.013633843                waigbacc=4.0293511e-011 aigc=0.010857174                laigc=-1.0328694e-011            waigc=3.6579227e-011 paigc=-4.4510785e-019            aigsd=0.0097493203               laigsd=-8.4558264e-012 waigsd=8.9138427e-011             paigsd=-7.2417184e-018            bigsd=0.00040255965 wbigsd=7.2174135e-011             tvoff=0.00222796                 ltvoff=-2.48268e-011 wtvoff=-3.84845e-010              ptvoff=7.77471e-018               kt1=-0.16439788 lkt1=-2.6158535e-009            wkt1=-2.1246722e-008            pkt1=1.836188e-015 kt2=-0.074660046               wkt2=1.2073887e-008             ua1=1.244775e-009 lua1=-9.5661544e-017            wua1=3.3386927e-016             pua1=-3.9031288e-023 ub1=-1.3102874e-018            wub1=-3.1450319e-025            uc1=5.2633566e-011 luc1=-3.2474182e-018            wuc1=-1.5426659e-017            puc1=8.3957862e-024 at=91460.738                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=2.2233406e-010 pcit=-7.8885408e-017            lu0=-5.0277018e-011            pu0=3.2067239e-018 lub=-3.7441797e-026            pub=-6.1802315e-033            laigbacc=-9.3054585e-011 paigbacc=1.8365782e-017             lbigsd=8.7083905e-012             pbigsd=-6.2069756e-018 lkt2=2.1092452e-009             pkt2=-1.6951909e-015            lub1=9.7326205e-026 pub1=4.179972e-032              lat=-0.0020203343              lvsat=0.0001432645 pvsat=1.2717605e-009             wat=-0.027609426               pat=2.506295e-009 letab=-7.4440366e-015            petab=6.573784e-020              leta0=0 peta0=0                          vsat_ss=2730.16                    vsat_ff=-3412.69 vsat_sf=1365.08                    vsat_fs=-1706.35                   wvsat_ss=9e-10 wvsat_ff=-3.6e-09                   wvsat_sf=-4.6e-09                   wvsat_fs=3.2e-09 ags_ss=0.100952                   ags_ff=-0.134603                  ags_sf=0.0504762 ags_fs=-0.0673016                 lags_ss=-8.6819e-09                lags_ff=1.15759e-08 lags_sf=-4.34096e-09               lags_fs=5.78794e-09                wags_ss=-4.7e-13 wags_ff=-4e-14                     wags_sf=-3.4e-14                   wags_fs=-2.2e-14 pags_ss=4.2e-21                    pags_ff=-3.2e-20                   pags_sf=-2.9e-21 pags_fs=3.9e-21                    lvsat_ss=-0.000578794               lvsat_ff=0.000723492 lvsat_sf=-0.000289396               lvsat_fs=0.000361746                pvsat_ss=-3.9e-16 pvsat_ff=4.8e-16                    pvsat_sf=-1.9e-16                   pvsat_fs=2.4e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.5 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.33161094 lvth0=1.508739e-009              wvth0=-2.3395704e-008            pvth0=8.5650313e-016 k2=0.0028869776               lk2=-1.0806248e-009            wk2=-2.038663e-008 pk2=2.0956602e-016             minv=-0.42453                   cit=0.0017617441 wcit=7.4504941e-010             voff=-0.18404726                lvoff=-1.6322619e-009 wvoff=-5.3322272e-009            pvoff=-2.9499557e-016            eta0=0.0096711111 weta0=-6.0440267e-009            etab=-0.033331574               wetab=-2.0487797e-008 u0=0.020071197                wu0=9.3234708e-010             ua=-1.8577834e-009 lua=2.1918621e-017             wua=-1.5800825e-017            pua=3.692403e-024 ub=1.8482499e-018             wub=5.8890086e-026             uc=9.0361317e-011 luc=3.7408231e-019             wuc=-2.126602e-017             puc=-3.3689852e-024 vsat=92997.42                   wvsat=-0.0097142557              a0=0.15508934 la0=-1.8326373e-007            wa0=2.8983906e-007             pa0=-7.7450564e-014 ags=2.9418746                  lags=-4.2630253e-009            wags=2.4394363e-008 pags=3.8623009e-015             keta=-0.25325657                lketa=1.3267172e-009 wketa=8.4490456e-008             pketa=-1.2020058e-015            pclm=1.1774384 lpclm=-7.2368549e-009            wpclm=8.4867508e-008             ppclm=-2.1007428e-015 pdiblc2=0.0008314353               lpdiblc2=2.9392181e-012             wpdiblc2=1.5167529e-009 ppdiblc2=-2.6470598e-017            aigbacc=0.012707239                waigbacc=4.3013323e-010 aigc=0.010880004                laigc=-1.2292098e-011            waigc=3.5710342e-011 paigc=-3.7038383e-019            aigsd=0.0097165306               laigsd=-5.6359142e-012 waigsd=-5.8997915e-011            paigsd=5.498007e-018              bigsd=0.00057383578 wbigsd=-6.3434298e-011            tvoff=0.00236881                 ltvoff=-3.69398e-011 wtvoff=-5.18913e-010              ptvoff=1.93045e-017               kt1=-0.14576412 lkt1=-4.2183569e-009            wkt1=-1.7318533e-008            pkt1=1.4983638e-015 kt2=-0.044516348               wkt2=-7.846098e-009             ua1=-1.4389381e-010 lua1=2.3763974e-017             wua1=-4.3726414e-017            pua1=-6.5580588e-024 ub1=2.4553188e-019             wub1=1.1217779e-025             uc1=6.4039967e-011 luc1=-4.2283687e-018            wuc1=3.9666723e-017             puc1=3.6577554e-024 at=54694.722                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.8958528e-010 pcit=-5.6502695e-017            lu0=-1.6153737e-010            pu0=-2.4304822e-017 lub=-2.3402892e-026            pub=-1.2982625e-032            laigbacc=-1.336663e-011 paigbacc=-1.5160434e-017            lbigsd=-6.0213572e-012            pbigsd=5.4553497e-018 lkt2=-4.8311287e-010            pkt2=1.7927814e-017             lub1=-3.647425e-026 pub1=5.1051552e-033             lat=0.001141543                lvsat=0.0020735622 pvsat=7.2497314e-010             wat=0.00044900751              pat=9.3269682e-011 letab=-1.0465637e-010            petab=9.414918e-016              leta0=0 peta0=0                          vsat_ss=-8166.62                   vsat_ff=9166.66 vsat_sf=-6166.67                   vsat_fs=7361.11                    wvsat_ss=-3.3e-09 wvsat_ff=-3.4e-09                   wvsat_sf=3.3e-09                    wvsat_fs=-3.3e-09 uc1_ss=3.08809e-11                luc1_ss=-2.65576e-18               wuc1_ss=-2.79781e-17 puc1_ss=2.40612e-24                lvsat_ss=0.000358334                lvsat_ff=-0.000358333 lvsat_sf=0.000358333                lvsat_fs=-0.000418055               pvsat_ss=2e-17 pvsat_ff=-5e-17                     pvsat_sf=-2e-17                     pvsat_fs=2e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.6 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.30220361 lvth0=2.9791054e-009             wvth0=-9.1689759e-009            pvth0=1.4516675e-016 k2=0.0243445                  lk2=-2.1535009e-009            wk2=-2.006168e-008 pk2=1.9331856e-016             minv=-0.42453                   cit=-0.0045157112 wcit=-2.2484899e-010            voff=-0.14249227                lvoff=-3.7100112e-009 wvoff=-2.3543495e-008            pvoff=6.1556781e-016             eta0=0.0063894239 weta0=-1.7516485e-008            etab=-0.066606929               wetab=-3.6208207e-009 u0=0.019207962                wu0=2.5351334e-010             ua=-1.8573846e-009 lua=2.1898681e-017             wua=1.3395283e-016             pua=-3.7952796e-024 ub=1.9751314e-018             wub=-3.8523954e-025            uc=1.363256e-010 luc=-1.9241317e-018            wuc=-1.0700166e-016            puc=9.1779664e-025 vsat=118207.52                  wvsat=0.015022329                a0=25.143416 la0=-1.43268e-006              wa0=-6.9954012e-006            pa0=2.8681145e-013 ags=2.8566141                  lags=0                          wags=1.0164038e-007 pags=0                          keta=0.38583123                 lketa=-3.0627673e-008 wketa=-1.230631e-007             pketa=9.1756719e-015             pclm=1.2544838 lpclm=-1.1089126e-008            wpclm=-4.1765732e-007            ppclm=2.3025499e-014 pdiblc2=0.00090041061              lpdiblc2=-5.0954733e-013            wpdiblc2=8.9556132e-010 ppdiblc2=4.5889832e-018             aigbacc=0.014157351                waigbacc=1.2692456e-010 aigc=0.010908688                laigc=-1.3726286e-011            waigc=1.0546504e-010 paigc=-3.8581188e-018            aigsd=0.0095556497               laigsd=2.4081327e-012 waigsd=-6.6520457e-012            paigsd=2.8807136e-018             bigsd=0.00071101376 wbigsd=-5.8425591e-013            tvoff=0.00170911                 ltvoff=-3.95461e-012 wtvoff=-3.17544e-010              ptvoff=9.23608e-018               kt1=-0.12942715 lkt1=-5.0352053e-009            wkt1=-2.1508872e-008            pkt1=1.7078807e-015 kt2=-0.040446264               wkt2=-5.2481179e-009            ua1=-6.4395344e-010 lua1=4.8766956e-017             wua1=1.2408111e-016             pua1=-1.4948435e-023 ub1=1.0234834e-018             wub1=-3.0943523e-025            uc1=-1.9059911e-011 luc1=-7.3374815e-020            wuc1=9.960556e-017              puc1=6.6081358e-025 at=51790.221                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=5.0345805e-010 pcit=-8.0077757e-018            lu0=-1.1837561e-010            pu0=9.6368647e-018 lub=-2.9746968e-026            pub=9.2238562e-033             laigbacc=-8.5872222e-011 paigbacc=-1.0959341e-030            lbigsd=-1.2880256e-011            pbigsd=2.3128475e-018 lkt2=-6.8661705e-010            pkt2=-1.1197119e-016            lub1=-7.5371828e-026 pub1=2.6185806e-032             lat=0.0012867681               lvsat=0.00081305723 pvsat=-5.118561e-010             wat=0.038343276                pat=-1.8014437e-009 letab=1.5591114e-009             petab=9.8142978e-017             leta0=1.6408436e-010 peta0=5.736229e-016              vsat_ss=-1000.01                   vsat_ff=6555.58 vsat_sf=1000.01                    vsat_fs=-1000.01                   wvsat_ss=4e-09 wvsat_ff=-5.4e-08                   wvsat_sf=-4e-09                     wvsat_fs=4e-09 uc1_ss=6.36147e-10                uc1_sf=6.58382e-10                luc1_ss=-3.29191e-17 luc1_sf=-3.29191e-17               wuc1_ss=-5.76349e-16               wuc1_sf=-5.96494e-16 puc1_ss=2.98247e-23                puc1_sf=2.98247e-23                at_ss=-30386.8 at_sf=-32919.1                   lat_ss=0.00151934                 lat_sf=0.00164595 lvsat_ss=2.52e-10                   lvsat_ff=-0.000227777               lvsat_sf=-2.52e-10 lvsat_fs=2.52e-10                   pvsat_ss=-7e-16                     pvsat_ff=-3e-16 pvsat_sf=7e-16                      pvsat_fs=-7e-16                     wat_ss=0.0275305 wat_sf=0.0298247                  pat_ss=-1.37652e-09               pat_sf=-1.49123e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.7 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.51415661 lvth0=-5.7109674e-009            wvth0=-1.9131231e-008            pvth0=5.5361919e-016 k2=0.058632005                lk2=-3.5592886e-009            wk2=-5.6075853e-008 pk2=1.6698996e-015             minv=-1.2228589                 cit=0.00336821 wcit=-1.9140649e-009            voff=-0.16530185                lvoff=-2.7748186e-009 wvoff=-2.7399391e-008            pvoff=7.7365954e-016             eta0=-0.033744288 weta0=6.502925e-009              etab=-0.054840027               wetab=-4.5790906e-009 u0=0.014721476                wu0=-2.7527587e-009            ua=-1.7671986e-009 lua=1.8201054e-017             wua=-8.6681642e-016            pua=3.7236259e-023 ub=1.0753454e-018             wub=9.2550837e-025             uc=1.5264757e-010 luc=-2.5933327e-018            wuc=-1.419227e-016             puc=2.3495594e-024 vsat=103593.2                   wvsat=0.0047850293               a0=-9.0888889 la0=-2.9155556e-008            ags=2.811264                   lags=1.8593547e-009 wags=1.4272759e-007             pags=-1.6845753e-015            keta=-1.0687934 lketa=2.9011937e-008             wketa=7.096135e-007              pketa=-2.4964069e-014 pclm=0.33141049                 lpclm=2.6756879e-008             wpclm=-3.8294956e-007 ppclm=2.1602481e-014             pdiblc2=-0.024899653               lpdiblc2=1.0572931e-009 wpdiblc2=2.2760419e-008             ppdiblc2=-8.9187019e-016            aigbacc=0.012212838 waigbacc=-1.2233558e-009            aigc=0.010233076                laigc=1.3973806e-011 waigc=4.1298185e-011             paigc=-1.2272777e-018            aigsd=0.0096650258 laigsd=-2.0762872e-012            waigsd=-3.154847e-010             paigsd=1.5542852e-017 bigsd=0.00053451097              wbigsd=-3.7723009e-010            tvoff=0.0025222 ltvoff=-3.72914e-011              wtvoff=-1.40745e-009              ptvoff=5.39221e-017 kt1=-0.18326523                lkt1=-2.8278443e-009            wkt1=1.7038951e-008 pkt1=1.2741998e-016             kt2=-0.070272464               wkt2=-1.4780667e-008 ua1=1.6419014e-009             lua1=-4.4953092e-017            wua1=-2.1386094e-016 pua1=-1.092811e-024             ub1=-1.632772e-018             wub1=2.6468257e-025 uc1=-9.1610048e-011            luc1=2.9011808e-018             wuc1=2.4065076e-016 puc1=-5.1220395e-024            at=87344.854                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.8021728e-010 pcit=6.1250077e-017             lu0=6.5570307e-011             pu0=1.3289402e-016 lub=7.1442611e-027             pub=-4.4516808e-032            laigbacc=-6.1471789e-012 paigbacc=5.5361493e-017             lbigsd=-5.643642e-012             pbigsd=1.7755327e-017 lkt2=5.3625716e-010             pkt2=2.7886333e-016             lub1=3.3534645e-026 pub1=2.6469762e-033             lat=-0.0001709719              lvsat=0.0014122442 pvsat=-9.2126812e-011            wat=-0.0055575362              pat=-1.5104436e-012 letab=1.0766684e-009             petab=1.3743204e-016             leta0=1.8095666e-009 peta0=-4.111729e-016             lminv=3.2731484e-008             vth0_ff=0.000595808 lvth0_ff=-2.44281e-11               wvth0_ff=-5.3718e-09                pvth0_ff=2.20244e-16 voff_ss=-0.00079441                voff_ff=0.00395276                 voff_mc=0.000993013 lvoff_ss=3.25708e-11                lvoff_ff=-1.62063e-10               lvoff_mc=-4.07135e-11 wvoff_ss=7.1624e-09                 wvoff_ff=-3.5812e-09                wvoff_mc=-8.953e-09 pvoff_ss=-2.93658e-16               pvoff_ff=1.46829e-16                pvoff_mc=3.67073e-16 eta0_sf=0.00790552                 eta0_fs=-0.00790552                weta0_sf=-7.1624e-09 weta0_fs=7.1624e-09                 u0_ss=3.97205e-05                u0_ff=-7.9441e-05 wu0_ss=-3.5812e-10                wu0_ff=7.1624e-10                 vsat_ss=-4555.55 vsat_ff=4754.16                    vsat_sf=4158.34                    vsat_fs=-4555.55 vsat_mc=-794.41                    wvsat_ss=-4e-09                     wvsat_ff=-0.0017906 wvsat_sf=0.00358121                 wvsat_fs=-4e-09                     wvsat_mc=0.0071624 uc1_ss=-7.59671e-10               uc1_sf=-6.58382e-10               luc1_ss=2.43095e-17 luc1_sf=2.10682e-17                wuc1_ss=6.88262e-16                wuc1_sf=5.96494e-16 puc1_ss=-2.20244e-23               puc1_sf=-1.90878e-23               at_ss=30386.8 at_sf=32919.1                    lu0_ss=-1.62854e-12               lu0_ff=3.25708e-12 pu0_ss=1.46829e-17                pu0_ff=-2.93658e-17               lat_ss=-0.000972379 lat_sf=-0.00105341                lvsat_ss=0.000145778                lvsat_ff=-0.000153921 lvsat_sf=-0.000129493               lvsat_fs=0.000145778                lvsat_mc=3.25708e-05 pvsat_ss=2.5e-16                    pvsat_ff=7.34147e-11                pvsat_sf=-1.4683e-10 pvsat_fs=2.5e-16                    pvsat_mc=-2.93658e-10               wat_ss=-0.0275305 wat_sf=-0.0298247                 pat_ss=8.80975e-10                pat_sf=9.5439e-10 leta0_sf=-3.24126e-10               leta0_fs=3.24126e-10                peta0_sf=2.93658e-16 peta0_fs=-2.93658e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_mac.8 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=0.36633405 lvth0=2.5496622e-012             wvth0=-1.4372961e-008            pvth0=-1.122623e-018 k2=-0.011424455               lk2=1.9359427e-013             wk2=-9.3630819e-009 pk2=-3.1955785e-019            minv=-0.42453                   cit=0.001 wcit=0                          voff=-0.15356225                lvoff=-2.8198957e-008 wvoff=2.3600819e-009             pvoff=4.3862699e-016             eta0=-3.3333333e-005 weta0=2.7482e-009                etab=-0.039217083               wetab=-5.3108965e-009 u0=0.0182607                  wu0=5.194098e-010              ua=-1.3897844e-009 lua=-2.8296734e-017            wua=-8.8112363e-017            pua=-1.7888129e-024 ub=1.74468e-018               wub=1.2531792e-025             uc=1.9787006e-010 luc=-6.7800372e-017            wuc=-2.8697994e-017            puc=1.0939079e-023 vsat=97416.667                  wvsat=0.0068705                  a0=1.9064821 la0=6.2437873e-007             wa0=3.5652724e-007             pa0=-5.6568713e-013 ags=0.97767742                 lags=1.5116977e-006             wags=1.1461206e-007 pags=-3.124878e-013             keta=-0.0054629007              lketa=-1.3377441e-007 wketa=2.4031314e-008             pketa=3.1042372e-014             pclm=0.22113952 lpclm=-4.0136228e-014            wpclm=1.620476e-007              ppclm=2.7347698e-020 pdiblc2=0.00030549794              lpdiblc2=1.7497405e-009             wpdiblc2=7.5999605e-011 ppdiblc2=-6.8369245e-016            aigbacc=0.013083                   aigc=0.010887774 laigc=-2.7738867e-011            waigc=2.1181202e-011             paigc=-6.3673645e-018 aigsd=0.0098232922               laigsd=2.1804743e-010             waigsd=-1.0042591e-010 paigsd=-1.3325048e-016            bigsd=0.00065466967              wbigsd=-1.4013072e-010 tvoff=0.00245242                 ltvoff=-2.41374e-010              wtvoff=-1.07532e-010 ptvoff=1.05836e-017               kt1=-0.16301745                lkt1=-1.8466811e-011 wkt1=1.1940762e-009             pkt1=1.2511572e-017             kt2=-0.058196667 wkt2=-1.09928e-009              ua1=1.6165237e-009             lua1=1.1672483e-017 wua1=-7.4829169e-017            pua1=-4.457858e-023             ub1=-1.5100267e-018 wub1=1.6709056e-025             uc1=1.0531266e-010             luc1=-1.1808675e-017 wuc1=1.2159937e-018             puc1=-1.0939079e-023            at=130000 jtsswgs='4.52e-005*(1+1.57*iboffn_flag)'                                   jtsswgd='4.52e-005*(1+1.57*iboffn_flag)' lcit=0                          pcit=0                          lu0=0 pu0=0                          lat=0                          lvsat=0 pvsat=0                          wat=0                          pat=0 leta0=0                          peta0=0                          vth0_mcl=-0.00223862 lvth0_mcl=-2.50406e-09               wvth0_mcl=1.22229e-09                pvth0_mcl=1.36721e-15 u0_mcl=-8.38413e-05               wu0_mcl=4.57774e-11                a0_sf=0.0139022 la0_sf=-1.25203e-07               wa0_sf=-7.59059e-09               pa0_sf=6.83608e-14 ags_ff=-0.252634                  lags_ff=2.2636e-07                 wags_ff=2.28887e-07 pags_ff=-2.05083e-13               lu0_mcl=7.51218e-11                pu0_mcl=-4.10165e-17 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.9 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.37435268 lvth0=-7.1821415e-009            wvth0=-1.9469834e-008            pvth0=4.5656751e-015 k2=-0.0016722338              lk2=-8.7377965e-009            wk2=-1.5220769e-008 pk2=5.2481678e-015             minv=-0.42453                   cit=-0.00012945866 wcit=-2.3383579e-010            voff=-0.19313222                lvoff=7.255735e-009 wvoff=1.1175343e-008             pvoff=-7.4598474e-015            eta0=-3.3333333e-005 weta0=2.7482e-009                etab=-0.039217083               wetab=-5.3108965e-009 u0=0.018054103                wu0=5.9703729e-010             ua=-1.2771924e-009 lua=-1.2917914e-016            wua=-1.2085188e-016            pua=2.7545794e-023 ub=1.5924536e-018             wub=2.4312104e-025             uc=1.4215437e-010 luc=-1.7879116e-017            wuc=-2.7384286e-017            puc=9.7619973e-024 vsat=97416.667                  wvsat=0.0068705                  a0=4.1990222 la0=-1.4297372e-006            wa0=-1.0919515e-006            pa0=7.3214979e-013 ags=3.4500608                  lags=-7.0355784e-007            wags=-1.1402811e-006 pags=8.1189649e-013             keta=-0.26921003                lketa=1.0254302e-007 wketa=1.3542589e-007             pketa=-6.8767169e-014            pclm=-0.21894081 lpclm=3.9431193e-007             wpclm=3.3627369e-007             ppclm=-1.5610655e-013 pdiblc2=0.0032114518               lpdiblc2=-8.5399419e-010            wpdiblc2=-1.64037e-009 ppdiblc2=8.5417476e-016             aigbacc=0.01315654                 waigbacc=-1.7976892e-010 aigc=0.010855405                laigc=1.2633608e-012             waigc=2.5886132e-011 paigc=-1.0582981e-017            aigsd=0.010412787                laigsd=-3.1013998e-010 waigsd=-5.0719654e-010            paigsd=2.31216e-016               bigsd=0.00080763314 wbigsd=-2.6931644e-010            tvoff=0.0022985                  ltvoff=-1.03459e-010 wtvoff=-9.43034e-011              ptvoff=-1.26906e-018              kt1=-0.16057455 lkt1=-2.2073028e-009            wkt1=9.6395062e-009             pkt1=-7.5545937e-015 kt2=-0.05620123                wkt2=-2.1887886e-009            ua1=2.1624338e-009 lua1=-4.7746295e-016            wua1=-2.9975416e-016            pua1=1.5695421e-022 ub1=-1.8685628e-018            wub1=3.1431041e-025             uc1=8.8036741e-011 luc1=3.670547e-018              wuc1=-9.7713778e-020            puc1=-9.7619973e-024 at=139911.11                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.011995e-009 pcit=2.0951687e-016             lu0=1.8511101e-010             pu0=-6.955423e-017 lub=1.3639486e-025             pub=-1.0555159e-031            laigbacc=-6.5892238e-011 paigbacc=1.6107295e-016             lbigsd=-1.3705527e-010            pbigsd=1.157504e-016 lkt2=-1.7879116e-009            pkt2=9.7619973e-016             lub1=3.2124834e-025 pub1=-1.3190899e-031            lat=-0.0088803556              lvsat=0 pvsat=0                          wat=0                          pat=0 leta0=0                          peta0=0                          vth0_mcl=-0.0100219 lvth0_mcl=4.46978e-09                wvth0_mcl=5.47197e-09                pvth0_mcl=-2.4405e-15 a0_sf=-0.250548                  la0_sf=1.11744e-07                wa0_sf=1.36799e-07 pa0_sf=-6.10125e-14               ags_ss=-0.0792892                 ags_ff=0.118934 ags_sf=-0.0495557                 ags_fs=0.0594669                  lags_ss=7.10427e-08 lags_ff=-1.06565e-07               lags_sf=4.44013e-08                lags_fs=-5.32818e-08 wags_ss=1.4e-13                    wags_ff=2.9e-13                    wags_sf=1.1e-14 wags_fs=4.7e-14                    pags_ss=-2.7e-20                   pags_ff=4e-20 pags_sf=-1.7e-20                   pags_fs=2.1e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.10 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.35677033 lvth0=6.5958816e-010             wvth0=-4.112038e-009             pvth0=-2.2839018e-015 k2=-0.019698093               lk2=-6.9826331e-010            wk2=-3.5513324e-009 pk2=4.3599242e-017             minv=-0.42453                   cit=0.00082639178 wcit=8.2763922e-010             voff=-0.15733177                lvoff=-8.7112619e-009 wvoff=-1.4953198e-008            pvoff=4.1934822e-015             eta0=-3.3333333e-005 weta0=2.7482e-009                etab=-0.039217083               wetab=-5.3108965e-009 u0=0.018333615                wu0=3.3651357e-010             ua=-1.4425706e-009 lua=-5.542046e-017             wua=-1.029386e-016             pua=1.9556473e-023 ub=1.9849999e-018             wub=3.0485054e-026             uc=1.2743419e-010 luc=-1.1313914e-017            wuc=-5.4964e-018               vsat=97416.667 wvsat=0.0068705                  a0=1.278416                   la0=-1.2714685e-007 wa0=9.4801156e-007             pa0=-1.7767371e-013            ags=1.3566288 lags=2.3011282e-007             wags=1.0024878e-006             pags=-1.4377844e-013 keta=0.033879061                lketa=-3.2634717e-008            wketa=-6.0091636e-008 pketa=1.8433648e-014             pclm=0.24901852                 lpclm=1.8560207e-007 wpclm=-6.3537444e-008            ppclm=2.2209214e-014             pdiblc2=0.0015745014 lpdiblc2=-1.239143e-010             wpdiblc2=-2.2314444e-010            ppdiblc2=2.2209214e-016 aigbacc=0.012367002                waigbacc=6.5942707e-010             aigc=0.010891989 laigc=-1.5052936e-011            waigc=-1.6840118e-011            paigc=8.4729263e-018 aigsd=0.0095200482               laigsd=8.8021574e-011             waigsd=1.5693372e-010 paigsd=-6.4986093e-017            bigsd=0.00047798077              wbigsd=9.2750076e-012 tvoff=0.00262691                 ltvoff=-2.49931e-010              wtvoff=-4.13819e-010 ptvoff=1.41235e-016               kt1=-0.14453695                lkt1=-9.3600729e-009 wkt1=-1.2319619e-008            pkt1=2.2391763e-015             kt2=-0.059917322 wkt2=-2.6516607e-010            ua1=1.2337578e-009             lua1=-6.3273492e-017 wua1=8.0095476e-017             pua1=-1.2458727e-023            ub1=-1.3055961e-018 wub1=4.0348744e-026             uc1=1.1450712e-010             luc1=-8.1352433e-018 wuc1=-3.1944889e-017            puc1=4.4418428e-024             at=166521.93 jtsswgs='4.52e-005*(1+1.57*iboffn_flag)'                                   jtsswgd='4.52e-005*(1+1.57*iboffn_flag)' lcit=5.8568566e-010             pcit=-2.6390099e-016            lu0=6.0448629e-011 pu0=4.663935e-017              lub=-3.8680792e-026            pub=-1.0715946e-032 laigbacc=2.8624204e-010             paigbacc=-2.1320846e-016            lbigsd=9.9696872e-012 pbigsd=-8.5013807e-018            lkt2=-1.3053429e-010            pkt2=1.1826407e-016 lub1=7.0165194e-026             pub1=-9.7220835e-033            lat=-0.020748782 lvsat=0                          pvsat=0                          wat=0.0034020673 pat=-1.517322e-009             leta0=0                          peta0=0 ags_ss=0.0981201                  ags_ff=-0.156239                  ags_sf=0.0681192 ags_fs=-0.0781196                 lags_ss=-8.08132e-09               lags_ff=1.61632e-08 lags_sf=-8.08131e-09               lags_fs=8.08138e-09                wags_ss=2.33e-13 wags_ff=-4.11e-13                  wags_sf=-4.33e-13                  wags_fs=7.44e-13 pags_ss=2.1e-20                    pags_ff=-2.8e-20                   pags_sf=1.1e-20 pags_fs=-1.4e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.11 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.36793845 lvth0=-1.7080546e-009            wvth0=-1.6540055e-008            pvth0=3.5083788e-016 k2=-0.021205586               lk2=-3.7867482e-010            wk2=-3.2287986e-009 pk2=-2.4777927e-017            minv=-0.42453                   cit=0.0031026765 wcit=-5.5457585e-010            voff=-0.18775889                lvoff=-2.2607141e-009 wvoff=7.2888759e-009             pvoff=-5.2183752e-016            eta0=-3.3333333e-005 weta0=2.7482e-009                etab=-0.039218146               wetab=-5.3102118e-009 u0=0.018846457                wu0=5.4994536e-010             ua=-1.7912587e-009 lua=1.8501423e-017             wua=-1.9941968e-017            pua=1.9611864e-024 ub=1.9621609e-018             wub=2.4487334e-026             uc=9.4536032e-011 luc=-4.3395054e-018            wuc=6.9359333e-019             puc=-1.3122786e-024 vsat=87333.917                  wvsat=0.0093943479               a0=2.9605515 la0=-4.8375959e-007            wa0=1.759546e-007              pa0=-1.3997638e-014 ags=2.1521147                  lags=6.1469815e-008             wags=4.8260137e-007 pags=-3.3562519e-014            keta=-0.072092773               lketa=-1.0168688e-008 wketa=2.6434674e-008             pketa=9.007003e-017              pclm=1.1209735 lpclm=7.4760847e-010             wpclm=5.0601778e-008             ppclm=-1.9883009e-015 pdiblc2=0.00012271958              lpdiblc2=1.8386345e-010             wpdiblc2=1.4247018e-009 ppdiblc2=-1.2725126e-016            aigbacc=0.015493214                waigbacc=-1.644296e-009 aigc=0.010872414                laigc=-1.0902961e-011            waigc=2.2771904e-011 paigc=7.5177657e-020             aigsd=0.010072107                laigsd=-2.9014961e-011 waigsd=-2.0330661e-010            paigsd=1.1384858e-017             bigsd=0.00059162159 wbigsd=-9.911599e-011             tvoff=0.0013873                  ltvoff=1.28663e-011 wtvoff=3.76795e-010               ptvoff=-2.63752e-017              kt1=-0.18349022 lkt1=-1.1019802e-009            wkt1=-3.9490651e-009            pkt1=4.6461879e-016 kt2=-0.069326197               wkt2=7.2414198e-009             ua1=1.5736759e-009 lua1=-1.3533613e-016            wua1=3.5885033e-017             pua1=-3.0861128e-024 ub1=-1.6476494e-018            wub1=-8.8531653e-027            uc1=6.2116334e-011 luc1=2.9716038e-018             wuc1=-2.4018047e-017            puc1=2.7613523e-024 at=67420.018                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.0311329e-010 pcit=2.9128608e-017             lu0=-4.8273802e-011            pu0=1.3918106e-018 lub=-3.383893e-026             pub=-9.4444292e-033            laigbacc=-3.7651492e-010 paigbacc=2.7518084e-016             lbigsd=-1.4122168e-011            pbigsd=1.4477511e-017 lkt2=1.8641472e-009             pkt2=-1.4731321e-015            lub1=1.4268051e-025 pub1=7.0872114e-034             lat=0.00026082397              lvsat=0.0021375429 pvsat=-5.3505575e-010            wat=-0.0058285346              pat=4.3956559e-010 letab=2.2531954e-013             petab=-1.4514596e-019            leta0=0 peta0=0                          vsat_ss=2730.16                    vsat_ff=-3412.69 vsat_sf=1365.08                    vsat_fs=-1706.35                   wvsat_ss=1.1e-09 wvsat_ff=1.1e-09                    wvsat_sf=-4.4e-09                   wvsat_fs=-4.4e-09 ags_ss=0.100952                   ags_ff=-0.134603                  ags_sf=0.0504764 ags_fs=-0.0673019                 lags_ss=-8.68194e-09               lags_ff=1.15759e-08 lags_sf=-4.34092e-09               lags_fs=5.78793e-09                wags_ss=-3.3e-13 wags_ff=-2.2e-13                   wags_sf=3.3e-14                    wags_fs=-1.1e-14 pags_ss=-5e-21                     pags_ff=7e-21                      pags_sf=-2.7e-21 pags_fs=3.6e-21                    lvsat_ss=-0.000578793               lvsat_ff=0.000723494 lvsat_sf=-0.000289396               lvsat_fs=0.000361746                pvsat_ss=-3.6e-16 pvsat_ff=4.4e-16                    pvsat_sf=-1.8e-16                   pvsat_fs=2.2e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.12 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.31746449 lvth0=2.6327057e-009             wvth0=-1.0579026e-008            pvth0=-1.6181062e-016 k2=-0.019938561               lk2=-4.8763892e-010            wk2=2.9330862e-010 pk2=-3.2767914e-016            minv=-0.42453                   cit=0.0028826081 wcit=-2.7045342e-010            voff=-0.18820602                lvoff=-2.2222609e-009 wvoff=-1.5643926e-009            pvoff=2.3954357e-016             eta0=-0.0015078704 weta0=4.0841306e-009             etab=-0.041568737               wetab=-1.3024927e-008 u0=0.02078717                 wu0=2.8367531e-010             ua=-1.7423946e-009 lua=1.4299106e-017             wua=-1.203431e-016             pua=1.0595684e-023 ub=1.9629882e-018             wub=-4.5062846e-026            uc=1.2214611e-010 luc=-6.7139722e-018            wuc=-5.0063043e-017            puc=3.0527922e-024 vsat=72328.909                  wvsat=0.0090114157               a0=-3.7727452 la0=9.5303926e-008             wa0=3.8484571e-006             pa0=-3.2983286e-013 ags=2.86688                    lags=0                          wags=9.233952e-008 pags=0                          keta=-0.21139815                lketa=1.8115741e-009 wketa=4.6566722e-008             pketa=-1.6412861e-015            pclm=1.0301296 lpclm=8.5601852e-009             wpclm=2.1832922e-007             ppclm=-1.6412861e-014 pdiblc2=0.0031139074               lpdiblc2=-7.3378704e-011            wpdiblc2=-5.5116678e-010 ppdiblc2=4.2673439e-017             aigbacc=0.0077556194               waigbacc=4.9163008e-009 aigc=0.010862813                laigc=-1.007728e-011             waigc=5.1285702e-011 paigc=-2.377009e-018             aigsd=0.009746402                laigsd=-1.004302e-012 waigsd=-8.6061361e-011            paigsd=1.3017664e-018             bigsd=0.00038641294 wbigsd=1.063708e-010              tvoff=0.00168781                 ltvoff=-1.29774e-011 wtvoff=9.80765e-011               ptvoff=-2.40544e-018              kt1=-0.16075121 lkt1=-3.0575346e-009            wkt1=-3.7402278e-009            pkt1=4.4665878e-016 kt2=-0.024469118               wkt2=-2.6008889e-008            ua1=-4.4825123e-010 lua1=3.8549606e-017             wua1=2.3202141e-016             pua1=-1.9953841e-023 ub1=7.2811242e-019             wub1=-3.2504018e-025            uc1=8.6489126e-011 luc1=8.755437e-019              wuc1=1.9327785e-017             puc1=-9.6638926e-025 at=49311.192                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.2203918e-010 pcit=4.6940783e-018             lu0=-2.1517518e-010            pu0=2.4291034e-017 lub=-3.3910079e-026            pub=-3.4631137e-033            laigbacc=2.8891819e-010 paigbacc=-2.8903048e-016            lbigsd=3.525776e-012              pbigsd=-3.1943531e-018 lkt2=-1.9935616e-009            pkt2=1.3863944e-015             lub1=-6.1635011e-026 pub1=2.7900804e-032             lat=0.0018181831               lvsat=0.0034279736 pvsat=-5.0212358e-010            wat=0.0053264865               pat=-5.1976623e-010 letab=2.0237612e-010             petab=6.6332037e-016             leta0=1.2681019e-010 peta0=-1.1489003e-016            vsat_ss=-8166.59                   vsat_ff=9166.72 vsat_sf=-6166.72                   vsat_fs=7361.15                    wvsat_ss=-1.78e-08 wvsat_ff=-8.44e-08                  wvsat_sf=-2.2e-09                   wvsat_fs=2.2e-09 lvsat_ss=0.000358335                lvsat_ff=-0.000358334               lvsat_sf=0.000358334 lvsat_fs=-0.000418059               pvsat_ss=3.9e-16                    pvsat_ff=2.2e-16 pvsat_sf=-3.9e-16                   pvsat_fs=3.9e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.13 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.30880329 lvth0=3.0657658e-009             wvth0=-1.5148286e-008            pvth0=6.6652354e-017 k2=0.033542374                lk2=-3.1616857e-009            wk2=-2.8394954e-008 pk2=1.106734e-015              minv=-0.42453                   cit=-0.0056992249 wcit=8.4741443e-010             voff=-0.20106853                lvoff=-1.5791353e-009 wvoff=2.9526594e-008             pvoff=-1.3150057e-015            eta0=-0.034262037 weta0=1.9313739e-008             etab=-0.054083128               wetab=-1.4967384e-008 u0=0.020662857                wu0=-1.0646221e-009            ua=-1.9267663e-009 lua=2.3517689e-017             wua=1.9681259e-016             pua=-5.2621006e-024 ub=1.5857358e-018             wub=-3.2447081e-026            uc=6.0888889e-012 luc=-9.1111111e-019            wuc=1.09928e-017               puc=2.5322685e-039 vsat=255738.07                  wvsat=-0.10958035                a0=47.661455 la0=-2.4764061e-006            wa0=-2.7396745e-005            pa0=1.2324272e-012 ags=2.6181467                  lags=1.2436667e-008             wags=3.1769192e-007 pags=-1.126762e-014             keta=0.30392593                 lketa=-2.395463e-008 wketa=-4.8856889e-008            pketa=3.1298944e-015             pclm=1.055436 lpclm=7.2948667e-009             wpclm=-2.3732002e-007            ppclm=6.3696012e-015 pdiblc2=0.0027988889               lpdiblc2=-5.7627778e-011            wpdiblc2=-8.2446e-010 ppdiblc2=5.63381e-017               aigbacc=0.020461009                waigbacc=-5.5841897e-009 aigc=0.011068828                laigc=-2.0378028e-011            waigc=-3.962167e-011 paigc=2.1683596e-018             aigsd=0.0098873655               laigsd=-8.0524761e-012 waigsd=-3.0718654e-010            paigsd=1.2358025e-017             bigsd=0.00076312614 wbigsd=-4.7798068e-011            tvoff=0.00103656                 ltvoff=1.9585e-011 wtvoff=2.91783e-010               ptvoff=-1.20908e-017              kt1=-0.12765069 lkt1=-4.7125605e-009            wkt1=-2.3118343e-008            pkt1=1.4155646e-015 kt2=-0.04681657                wkt2=5.2337942e-010             ua1=-3.7917609e-010 lua1=3.5095849e-017             wua1=-1.1580717e-016            pua1=-2.5624122e-024 ub1=5.5540137e-019             wub1=1.1464712e-025             uc1=7.0981333e-011 luc1=1.6509333e-018             wuc1=1.8028192e-017             puc1=-9.014096e-025 at=145921.41                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=5.5113083e-010 pcit=-5.1199314e-017            lu0=-2.0895954e-010            pu0=9.1705907e-017 lub=-1.5047456e-026            pub=-4.0939019e-033            laigbacc=-3.463513e-010 paigbacc=2.3599404e-016             lbigsd=-1.5309884e-011            pbigsd=4.5140903e-018 lkt2=-8.7618898e-010            pkt2=5.9780984e-017             lub1=-5.2999459e-026 pub1=5.9164395e-033             lat=-0.0030123277              lvsat=-0.0057424846 pvsat=5.4274648e-009             wat=-0.046939578               pat=2.093537e-009 letab=8.2809567e-010             petab=7.6044322e-016             leta0=1.7645185e-009 peta0=-8.7637044e-016            vsat_ss=-1000.02                   vsat_ff=6555.61 vsat_sf=1000.02                    vsat_fs=-1000.02                   wvsat_ss=-1.1e-09 wvsat_ff=-1.89e-08                  wvsat_sf=1.1e-09                    wvsat_fs=-1.1e-09 lvsat_ss=-4e-11                     lvsat_ff=-0.000227776               lvsat_sf=4e-11 lvsat_fs=-4e-11                     pvsat_ss=5.6e-16                    pvsat_ff=4.4e-16 pvsat_sf=-5.6e-16                   pvsat_fs=5.6e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.14 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.61234364 lvth0=-9.3793883e-009            wvth0=-1.0808868e-007            pvth0=3.8772085e-015 k2=-0.019657981               lk2=-9.8047113e-010            wk2=1.4854875e-008 pk2=-6.6650899e-016            minv=-1.7066542                 cit=0.0035090097 wcit=-2.0416295e-009            voff=-0.21597915                lvoff=-9.6779975e-010 wvoff=1.8514247e-008             pvoff=-8.6349952e-016            eta0=-0.010270926 weta0=-1.4763941e-008            etab=-0.0747036                 wetab=1.3417307e-008 u0=0.006609187                wu0=4.5969752e-009             ua=-3.3649749e-009 lua=8.2484245e-017             wua=5.8076895e-016             pua=-2.1004312e-023 ub=2.409965e-018              wub=-2.8365699e-025            uc=5.437037e-012 luc=-8.8438518e-019            wuc=-8.5499556e-018            puc=8.0125298e-025 vsat=61677.321                  wvsat=0.042760818                a0=-22.47627 la0=3.9924063e-007             wa0=1.2128967e-005             pa0=-3.8812694e-013 ags=3.1156133                  lags=-7.9594667e-009            wags=-1.3301288e-007 pags=7.2112768e-015             keta=-0.15411111                lketa=-5.1751111e-009 wketa=-1.1908867e-007            pketa=6.0093973e-015             pclm=0.051230668 lpclm=4.8467285e-008             wpclm=-1.2910664e-007            ppclm=1.9328525e-015 pdiblc2=-0.0030807407              lpdiblc2=1.8343704e-010             wpdiblc2=2.9924844e-009 ppdiblc2=-1.0015662e-016            aigbacc=0.0046710167               waigbacc=5.6095342e-009 aigc=0.0099105511               laigc=2.7111305e-011             waigc=3.3350544e-010 paigc=-1.3129852e-017            aigsd=0.0085574674               laigsd=4.6473345e-011 waigsd=6.8796321e-010             paigsd=-2.8443115e-017            bigsd=-0.00073848122 wbigsd=7.7610084e-010             tvoff=-0.000394327               ltvoff=7.82514e-011 wtvoff=1.23493e-009               ptvoff=-5.07597e-017              kt1=-0.19377031 lkt1=-2.0016562e-009            wkt1=2.655656e-008              pkt1=-6.2110647e-016 kt2=-0.096549819               wkt2=9.0266156e-009             ua1=1.9311713e-009 lua1=-5.9628394e-017            wua1=-4.7593948e-016            pua1=1.2203013e-023 ub1=-1.7040285e-018            wub1=3.2924092e-025             uc1=2.1344593e-011 luc1=3.6860397e-018             wuc1=1.3831385e-016             puc1=-5.8331217e-024 at=104396.74                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.7359321e-010 pcit=6.7251486e-017             lu0=3.6724095e-010             pu0=-1.4041958e-016 lub=-4.8840852e-026            pub=6.2057043e-033             laigbacc=3.010384e-010 paigbacc=-2.2294864e-016            lbigsd=4.6256018e-011             pbigsd=-2.9265765e-017 lkt2=1.1628742e-009             pkt2=-2.888517e-016             lub1=3.9637165e-026 pub1=-2.8819067e-033            lat=-0.0013098164              lvsat=0.0022140062 pvsat=-8.1852318e-010            wat=-0.021006545               pat=1.0302826e-009 letab=1.673535e-009              petab=-4.0332912e-016            leta0=7.8088296e-010 peta0=5.2081444e-016             lminv=5.2567093e-008             wminv=4.3831857e-007 pminv=-1.7971062e-014            vth0_ss=0.00539259                 vth0_ff=-0.0215111 lvth0_ss=-2.21096e-10               lvth0_ff=8.81955e-10                wvth0_ss=-4.88569e-09 wvth0_ff=1.46571e-08                pvth0_ss=2.00313e-16                pvth0_ff=-6.0094e-16 voff_ss=0.00711112                 voff_ff=0.0161778                  voff_mc=-0.0223704 lvoff_ss=-2.91555e-10               lvoff_ff=-6.63289e-10               lvoff_mc=9.17185e-10 wvoff_ss=-2.2e-15                   wvoff_ff=-1.46571e-08               wvoff_mc=1.22142e-08 pvoff_ss=-4.9e-22                   pvoff_ff=6.0094e-16                 pvoff_mc=-5.00783e-16 u0_ss=-0.00197333                u0_ff=0.000980741                u0_sf=-0.000539259 wu0_ss=1.46571e-09                wu0_ff=-2.44285e-10               wu0_sf=4.88569e-10 vsat_ss=-9948.14                   vsat_ff=2777.78                    vsat_sf=2718.42 vsat_fs=-4555.54                   vsat_mc=4414.8                     wvsat_ss=0.00488571 wvsat_ff=-1.1e-09                   wvsat_sf=0.00488567                 wvsat_fs=1.1e-09 wvsat_mc=0.00244282                 lu0_ss=8.09067e-11                lu0_ff=-4.02104e-11 lu0_sf=2.21096e-11                pu0_ss=-6.00939e-17               pu0_ff=1.00156e-17 pu0_sf=-2.00313e-17               lvsat_ss=0.000366874                lvsat_ff=-7.28887e-05 lvsat_sf=-7.04594e-05               lvsat_fs=0.000145778                lvsat_mc=-0.000181007 pvsat_ss=-2.00313e-10               pvsat_ff=-2.4e-16                   pvsat_sf=-2.00313e-10 pvsat_fs=2.4e-16                    pvsat_mc=-1.00157e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.15 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.36928647 lvth0=-2.2255151e-013            wvth0=-1.5984982e-008            pvth0=3.9100567e-019 k2=-0.024559724               lk2=-2.8680044e-013            wk2=-2.1912251e-009 pk2=-5.7262336e-020            minv=-0.42453                   cit=0.0011022222 wcit=-5.5813333e-011            voff=-0.16400548                lvoff=-2.5956892e-008 wvoff=8.0620892e-009             pvoff=-7.8554039e-016            eta0=0.005 weta0=0                          etab=-0.0451168                 wetab=-2.0896512e-009 u0=0.018566978                wu0=3.5218213e-010             ua=-1.5673084e-009 lua=1.3970499e-017             wua=8.815736e-018              pua=-2.4866722e-023 ub=1.8928311e-018             wub=4.4427413e-026             uc=1.6256979e-010 luc=-5.5903242e-017            wuc=-9.4240469e-018            puc=4.4432463e-024 vsat=97733.333                  wvsat=0.0066976                  a0=1.9100608 la0=2.6177666e-007             wa0=3.5457327e-007             pa0=-3.677064e-013 ags=1.179271                   lags=1.1171887e-006             wags=4.5419901e-009 pags=-9.7085892e-014            keta=0.050458333                lketa=-9.208405e-008 wketa=-6.5016795e-009            pketa=8.279434e-015              pclm=0.58736953 lpclm=2.0123398e-014             wpclm=-3.7913991e-008            ppclm=-5.5540578e-021 pdiblc2=0.00060299698              lpdiblc2=-9.2656085e-010            wpdiblc2=-8.6434871e-011 ppdiblc2=7.775681e-016              aigbacc=0.0132118                  waigbacc=-7.03248e-011 aigc=0.010880211                laigc=-4.3994604e-011            waigc=2.5310644e-011 paigc=2.5082681e-018             aigsd=0.0096395746               laigsd=-1.0922171e-010 waigsd=-1.1606595e-013            paigsd=4.5438469e-017             bigsd=0.00037227022 wbigsd=1.4059379e-011             tvoff=0.00234906                 ltvoff=-4.13756e-010 wtvoff=-5.1099e-011               ptvoff=1.04704e-016               kt1=-0.1596657 lkt1=9.2698101e-012             wkt1=-6.3597936e-010            pkt1=-2.6326234e-018 kt2=-0.06021                   ua1=1.3921794e-009             lua1=-2.9933454e-017 wua1=4.7662789e-017             pua1=-2.1861738e-023            ub1=-1.07244e-018 wub1=-7.183176e-026             uc1=1.1115817e-010             luc1=-6.4394873e-017 wuc1=-1.9756542e-018            puc1=1.7772985e-023             at=130000 jtsswgs='4.52e-005*(1+1.57*iboffn_flag)'                                   jtsswgd='4.52e-005*(1+1.57*iboffn_flag)' lcit=0                          pcit=0                          lu0=0 pu0=0                          lat=0                          lvsat=0 pvsat=0                          wat=0                          pat=0 leta0=0                          peta0=0                          ags_ff=0.109814 lags_ff=-9.83936e-08               wags_ff=3.09898e-08                pags_ff=-2.77669e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.16 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.37737077 lvth0=-7.2437606e-009            wvth0=-2.1117714e-008            pvth0=4.5993192e-015 k2=-0.025721338               lk2=1.0405193e-009             wk2=-2.0899581e-009 pk2=-9.0792539e-017            minv=-0.42453                   cit=-0.00042683537 wcit=-7.1468105e-011            voff=-0.19810469                lvoff=4.5959936e-009 wvoff=1.3890313e-008             pvoff=-6.0076286e-015            eta0=0.005 weta0=0                          etab=-0.0451168                 wetab=-2.0896512e-009 u0=0.018501542                wu0=3.5273531e-010             ua=-1.4493836e-009 lua=-9.1690069e-017            wua=-2.6835472e-017            pua=7.0767601e-024 ub=1.8968903e-018             wub=7.6898618e-026             uc=1.0423032e-010 luc=-3.6310787e-018            wuc=-6.6777553e-018            puc=1.982569e-024 vsat=97733.333                  wvsat=0.0066976                  a0=2.0987062 la0=9.275038e-008              wa0=5.4821096e-008             pa0=-9.9128449e-014 ags=1.3731051                  lags=9.4351326e-007             wags=-6.2633256e-009 pags=-8.7404329e-014            keta=-0.023985688               lketa=-2.5382207e-008 wketa=1.5333982e-009             pketa=1.0800044e-015             pclm=0.44402472 lpclm=1.2843698e-007             wpclm=-2.5705488e-008            ppclm=-1.0938824e-014 pdiblc2=-0.00092005926             lpdiblc2=4.3809754e-010             wpdiblc2=6.1543502e-010 ppdiblc2=1.4869267e-016             aigbacc=0.012822359                waigbacc=2.6939236e-012 aigc=0.010833266                laigc=-1.9325844e-012            waigc=3.7973884e-011 paigc=-8.8379951e-018            aigsd=0.0092673005               laigsd=2.2433584e-010 waigsd=1.1823914e-010             paigsd=-6.0607793e-017            bigsd=0.00025395833 wbigsd=3.2990011e-011             tvoff=0.00183901                 ltvoff=4.32505e-011 wtvoff=1.56576e-010               ptvoff=-8.13722e-017              kt1=-0.14085543 lkt1=-1.6844728e-008            wkt1=-1.1271324e-009            pkt1=4.3744046e-016 kt2=-0.062035671               wkt2=9.9681621e-010             ua1=1.5423289e-009 lua1=-1.6446735e-016            wua1=3.8823115e-017             pua1=-1.394139e-023 ub1=-1.0978191e-018            wub1=-1.0651565e-025            uc1=5.2733377e-011 luc1=-1.2046261e-017            wuc1=1.9177923e-017             puc1=-1.1806198e-024 at=139911.11                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.3700356e-009 pcit=1.4026676e-017             lu0=5.8630081e-011             pu0=-4.9564225e-019 lub=-3.6369989e-027            pub=-2.90942e-032              laigbacc=3.4893877e-010 paigbacc=-6.5424776e-017            lbigsd=1.0600746e-010             pbigsd=-1.6961847e-017 lkt2=1.635801e-009              pkt2=-8.9314732e-016            lub1=2.2739631e-026 pub1=3.1076769e-032             lat=-0.0088803556              lvsat=0 pvsat=0                          wat=0                          pat=0 leta0=0                          peta0=0                          ags_ss=-0.0792891 ags_ff=0.118934                   ags_sf=-0.0495552                 ags_fs=0.0594669 lags_ss=7.10424e-08                lags_ff=-1.06565e-07               lags_sf=4.44018e-08 lags_fs=-5.32818e-08               wags_ss=2.8e-14                    wags_ff=-4.2e-14 wags_sf=-7e-15                     wags_fs=2.9e-14                    pags_ss=-2e-20 pags_ff=3.1e-20                    pags_sf=1.2e-20                    pags_fs=-3.5e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.17 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.371743 lvth0=-4.7337724e-009            wvth0=-1.2287118e-008            pvth0=6.6087314e-016 k2=-0.02163383                lk2=-7.8250915e-010            wk2=-2.49442e-009 pk2=8.9597472e-017             minv=-0.42453                   cit=0.0021809227 wcit=8.806533e-011              voff=-0.19086765                lvoff=1.3682756e-009 wvoff=3.3573904e-009             pvoff=-1.3099453e-015            eta0=0.005 weta0=0                          etab=-0.0451168                 wetab=-2.0896512e-009 u0=0.018418                   wu0=2.9043923e-010             ua=-1.5722961e-009 lua=-3.6871101e-017            wua=-3.2108484e-017            pua=9.4285237e-024 ub=1.9642724e-018             wub=4.1802279e-026             uc=1.2145641e-010 luc=-1.1313914e-017            wuc=-2.2325333e-018            vsat=97733.333 wvsat=0.0066976                  a0=3.8029478                  la0=-6.6734137e-007 wa0=-4.3038282e-007            pa0=1.172725e-013              ags=3.8653186 lags=-1.6801394e-007            wags=-3.6725683e-007            pags=7.3598775e-014 keta=-0.085450541               lketa=2.031117e-009              wketa=5.0623266e-009 pketa=-4.9389762e-016            pclm=0.40061159                 lpclm=1.4779923e-007 wpclm=-1.4630726e-007            ppclm=4.2849566e-014             pdiblc2=-0.0011276353 lpdiblc2=5.3067647e-010             wpdiblc2=1.2522222e-009             ppdiblc2=-1.3531442e-016 aigbacc=0.013493036                waigbacc=4.4612504e-011             aigc=0.010818943 laigc=4.4559044e-012             waigc=2.3043179e-011             paigc=-2.1789004e-018 aigsd=0.0098830087               laigsd=-5.027e-011                waigsd=-4.12427e-011 paigsd=1.0521106e-017             bigsd=0.00046590754              wbigsd=1.5866987e-011 tvoff=0.00181497                 ltvoff=5.39725e-011               wtvoff=2.95001e-011 ptvoff=-2.46965e-017              kt1=-0.16246614                lkt1=-7.2063538e-009 wkt1=-2.530283e-009             pkt1=1.0632457e-015             kt2=-0.063098898 wkt2=1.4719741e-009             ua1=1.228772e-009              lua1=-2.4620968e-017 wua1=8.2817766e-017             pua1=-3.3563005e-023            ub1=-9.6218916e-019 wub1=-1.4715142e-025            uc1=4.2747684e-011             luc1=-7.5926423e-018 wuc1=7.2357646e-018             puc1=4.1455827e-024             at=179350.21 jtsswgs='4.52e-005*(1+1.57*iboffn_flag)'                                   jtsswgd='4.52e-005*(1+1.57*iboffn_flag)' lcit=2.0697549e-010             pcit=-5.7125237e-017            lu0=9.5889915e-011 pu0=2.7288408e-017             lub=-3.3689425e-026            pub=-1.3441232e-032 laigbacc=4.9817141e-011             paigbacc=-8.4120463e-017            lbigsd=1.1478107e-011 pbigsd=-9.3249777e-018            lkt2=2.1100002e-009             pkt2=-1.1050677e-015 lub1=-3.77513e-026              pub1=4.9200322e-032             lat=-0.026470193 lvsat=0                          pvsat=0                          wat=-0.0036021715 pat=1.6065685e-009             leta0=0                          peta0=0 ags_ss=0.09812                    ags_ff=-0.15624                   ags_sf=0.0681196 ags_fs=-0.0781193                 lags_ss=-8.08136e-09               lags_ff=1.61627e-08 lags_sf=-8.08135e-09               lags_fs=8.08145e-09                wags_ss=4.4e-14 wags_ff=-5.9e-14                   wags_sf=2.2e-14                    wags_fs=-3e-14 pags_ss=-5.8e-20                   pags_ff=-2.2e-20                   pags_sf=9e-22 pags_fs=3.88e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.18 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.35768883 lvth0=-1.7542886e-009            wvth0=-1.0943762e-008            pvth0=3.7608164e-016 k2=-0.023765106               lk2=-3.3067854e-010            wk2=-1.8313003e-009 pk2=-5.0983899e-017            minv=-0.42453                   cit=0.0026571102 wcit=-3.1129665e-010            voff=-0.16652262                lvoff=-3.7928718e-009 wvoff=-4.3061277e-009            pvoff=3.1472056e-016             eta0=0.005 weta0=0                          etab=-0.045116274               wetab=-2.0898341e-009 u0=0.018811795                wu0=5.6887076e-010             ua=-1.8907356e-009 lua=3.0638066e-017             wua=3.4372384e-017             pua=-4.6654205e-024 ub=2.1016884e-018             wub=-5.1694664e-026            uc=9.7523033e-011 luc=-6.2400387e-018            wuc=-9.3730963e-019            puc=-2.7458742e-025 vsat=90337.555                  wvsat=0.0077543616               a0=2.9465697 la0=-4.8578923e-007            wa0=1.8358866e-007             pa0=-1.2889457e-014 ags=3.0579388                  lags=3.1505668e-009             wags=-1.1978604e-008 pags=-1.7202095e-015            keta=-0.032098394               lketa=-9.2795382e-009 wketa=4.5977429e-009             pketa=-3.9540589e-016            pclm=1.055612 lpclm=8.9391464e-009             wpclm=8.6289185e-008             ppclm=-6.4608806e-015 pdiblc2=0.0014262152               lpdiblc2=-1.0739838e-011            wpdiblc2=7.1299318e-010 ppdiblc2=-2.0997862e-017            aigbacc=0.012601331                waigbacc=-6.5328178e-011 aigc=0.010876904                laigc=-7.8319913e-012            waigc=2.0319929e-011 paigc=-1.6015715e-018            aigsd=0.0096683452               laigsd=-4.7613443e-012 waigsd=1.7147505e-011             paigsd=-1.857617e-018             bigsd=0.00042643954 wbigsd=-8.9265896e-012            tvoff=0.00240344                 ltvoff=-7.07819e-011 wtvoff=-1.78015e-010              ptvoff=1.92967e-017               kt1=-0.20314176 lkt1=1.4168791e-009             wkt1=6.7806796e-009             pkt1=-9.106784e-016 kt2=-0.047349712               wkt2=-4.7577412e-009            ua1=2.0877636e-009 lua1=-2.0672719e-016            wua1=-2.4480681e-016            pua1=3.5893406e-023 ub1=-2.2335539e-018            wub1=3.1105066e-025             uc1=-6.9653807e-011 luc1=1.6236474e-017             wuc1=4.7928451e-017             puc1=-4.4812668e-024 at=47300.39                   jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.0602374e-010 pcit=2.7539504e-017             lu0=1.2405477e-011             pu0=-3.1739076e-017 lub=-6.282162e-026             pub=6.3801196e-033             laigbacc=2.3885849e-010 paigbacc=-6.0813039e-017            lbigsd=1.9845323e-011             pbigsd=-4.0687395e-018 lkt2=-1.2288271e-009            pkt2=2.1563189e-016             lub1=2.3177802e-025 pub1=-4.7938519e-032            lat=0.0015243685               lvsat=0.001567905 pvsat=-2.2403346e-010            wat=0.0051567823               pat=-2.5032971e-010 letab=-1.1151424e-013            petab=3.8765284e-020             leta0=0 peta0=0                          vsat_ss=2730.16                    vsat_ff=-3412.69 vsat_sf=1365.08                    vsat_fs=-1706.35                   wvsat_ss=2.6e-09 wvsat_ff=-7e-10                     wvsat_sf=3e-10                      wvsat_fs=-3.7e-10 ags_ss=0.100952                   ags_ff=-0.134604                  ags_sf=0.0504761 ags_fs=-0.0673018                 lags_ss=-8.68186e-09               lags_ff=1.15759e-08 lags_sf=-4.34095e-09               lags_fs=5.78794e-09                wags_ss=-1.1e-14 wags_ff=-1.9e-14                   wags_sf=4.4e-14                    wags_fs=4.1e-14 pags_ss=-4e-22                     pags_ff=6e-22                      pags_sf=-2e-22 pags_fs=3e-22                      lvsat_ss=-0.000578794               lvsat_ff=0.00072349 lvsat_sf=-0.000289397               lvsat_fs=0.000361746                pvsat_ss=-3e-17 pvsat_ff=4e-17                      pvsat_sf=-1e-17                     pvsat_fs=-4.8e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.19 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.30725465 lvth0=2.5830509e-009             wvth0=-5.0044509e-009            pvth0=-1.346991e-016 k2=-0.014501214               lk2=-1.1273733e-009            wk2=-2.6754832e-009 pk2=2.1615833e-017             minv=-0.42453                   cit=0.00206425 wcit=1.7637013e-010             voff=-0.18960487                lvoff=-1.8077976e-009 wvoff=-8.0061637e-010            pvoff=1.3246586e-017             eta0=0.0055462963 weta0=2.3255556e-010             etab=-0.054012724               wetab=-6.2305101e-009 u0=0.022181631                wu0=-4.7770012e-010            ua=-1.9008624e-009 lua=3.1508972e-017             wua=-3.3819675e-017            pua=1.1990967e-024 ub=1.8808588e-018             wub=-2.2015259e-028            uc=1.4452099e-011 luc=9.0406173e-019             wuc=8.7378874e-018             puc=-1.1066544e-024 vsat=64722.138                  wvsat=0.013164713                a0=1.390438 la0=-3.519619e-007             wa0=1.0293591e-006             pa0=-8.5625715e-014 ags=3.0945733                  lags=0                          wags=-3.198104e-008 pags=0                          keta=-0.18290124                lketa=3.6895062e-009 wketa=3.1007407e-008             pketa=-2.666637e-015             pclm=1.3811605 lpclm=-1.9058025e-008            wpclm=2.666637e-008              ppclm=-1.3333185e-015 pdiblc2=0.00047911111              lpdiblc2=7.0711111e-011             wpdiblc2=8.87432e-010 ppdiblc2=-3.59996e-017              aigbacc=0.019624157                waigbacc=-1.5639206e-009 aigc=0.010961516                laigc=-1.5108583e-011            waigc=-2.6062811e-012 paigc=3.7008256e-019             aigsd=0.0095816993               laigsd=2.690208e-012 waigsd=3.866331e-012              paigsd=-7.1543605e-019            bigsd=0.00072046174 wbigsd=-7.601985e-011             tvoff=0.00192251                 ltvoff=-2.94225e-011 wtvoff=-3.00722e-011              ptvoff=6.57359e-018               kt1=-0.13401722 lkt1=-4.527832e-009             wkt1=-1.833699e-008             pkt1=1.2494412e-015 kt2=-0.065116363               wkt2=-3.8154925e-009            ua1=-9.9231676e-010 lua1=5.8159718e-017             wua1=5.2908119e-016             pua1=-3.0660962e-023 ub1=1.4405679e-018             wub1=-7.1404085e-025            uc1=2.0832166e-010 luc1=-7.6694163e-018            wuc1=-4.7192778e-017            puc1=3.6991589e-024 at=40943.097                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.5700972e-010 pcit=-1.439984e-017             lu0=-2.7740043e-010            pu0=5.8266019e-017 lub=-4.3830272e-026            pub=1.9533116e-033             laigbacc=-3.6510451e-010 paigbacc=6.806591e-017              lbigsd=-5.4405865e-012            pbigsd=1.7012808e-018 lkt2=2.9910481e-010             pkt2=1.345985e-016              lub1=-8.4196451e-026 pub1=4.0219351e-032             lat=0.0020710957               lvsat=0.0037708309 pvsat=-6.8932367e-010            wat=0.0098954661               pat=-6.5785652e-010 letab=7.6498318e-010             petab=3.5613691e-016             leta0=-4.6981482e-011 peta0=-1.9999778e-017            vsat_ss=-8166.75                   vsat_ff=9166.63 vsat_sf=-6166.7                    vsat_fs=7361.11                    wvsat_ss=-8.81e-09 wvsat_ff=-4e-10                     wvsat_sf=7.81e-09                   wvsat_fs=-8.81e-09 lvsat_ss=0.000358334                lvsat_ff=-0.000358338               lvsat_sf=0.000358332 lvsat_fs=-0.000418055               pvsat_ss=-2.26e-16                  pvsat_ff=-1.5e-16 pvsat_sf=-2.74e-16                  pvsat_fs=2.74e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.20 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.29293296 lvth0=3.2991354e-009             wvth0=-6.4830844e-009            pvth0=-6.0767427e-017 k2=-0.017750079               lk2=-9.6493004e-010            wk2=-3.8927496e-010 pk2=-9.269458e-017             minv=-0.42453                   cit=-0.0088343174 wcit=2.5591749e-009             voff=-0.11340058                lvoff=-5.6180124e-009 wvoff=-1.8340107e-008            pvoff=8.9022114e-016             eta0=0.01445679 weta0=-7.2867407e-009            etab=-0.10331552                wetab=1.1913503e-008 u0=0.012824773                wu0=3.214972e-009              ua=-1.0491228e-009 lua=-1.1078008e-017            wua=-2.8238075e-016            pua=1.362715e-023 ub=5.9876464e-019             wub=5.0643916e-025             uc=-4.2380247e-011 luc=3.745679e-018              wuc=3.7456948e-017             puc=-2.5426074e-024 vsat=52680.309                  wvsat=0.0012891869               a0=7.942269 la0=-6.7955345e-007            wa0=-5.7100693e-006            pa0=2.5134571e-013 ags=3.4262178                  lags=-1.6582222e-008            wags=-1.2351491e-007 pags=4.5766933e-015             keta=0.67444444                 lketa=-3.9177778e-008 wketa=-2.5116e-007               pketa=1.1441733e-014             pclm=0.50166395 lpclm=2.4916803e-008             wpclm=6.5039516e-008             ppclm=-3.2519758e-015 pdiblc2=0.0023792593               lpdiblc2=-2.4296296e-011            wpdiblc2=-5.9534222e-010 ppdiblc2=3.8139111e-017             aigbacc=0.013468548                waigbacc=-1.766306e-009 aigc=0.010993091                laigc=-1.6687362e-011            waigc=1.7302567e-012 paigc=1.5325566e-019             aigsd=0.0094942236               laigsd=7.0639903e-012 waigsd=-9.253108e-011             paigsd=4.1044345e-018             bigsd=0.0011014 wbigsd=-2.3249561e-010            tvoff=0.00188079                 ltvoff=-2.73362e-011 wtvoff=-1.69164e-010              ptvoff=1.35282e-017               kt1=-0.13297069 lkt1=-4.5801581e-009            wkt1=-2.0213623e-008            pkt1=1.3432728e-015 kt2=-0.023552543               wkt2=-1.2178779e-008            ua1=-5.0510946e-010 lua1=3.3799353e-017             wua1=-4.704755e-017             pua1=-1.8545254e-024 ub1=5.9100484e-019             wub1=9.5207624e-026             uc1=-5.682963e-011 luc1=5.5881482e-018             wuc1=8.7812978e-017             puc1=-3.0511289e-024 at=44272.245                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=7.0193809e-010 pcit=-1.3354008e-016            lu0=1.9044247e-010             pu0=-1.2636759e-016 lub=2.0274435e-026             pub=-2.3379654e-032            laigbacc=-5.7324074e-011 paigbacc=7.8185178e-017             lbigsd=-2.44875e-011              pbigsd=9.5250687e-018 lkt2=-1.7790862e-009            pkt2=5.5276285e-016             lub1=-4.17183e-026 pub1=-2.4307327e-034            lat=0.0019046383               lvsat=0.0043729223 pvsat=-9.5547373e-011            wat=0.0085608639               pat=-5.9112641e-010 letab=3.2301231e-009             petab=-5.5106375e-016            leta0=-4.9250617e-010 peta0=3.5596504e-016             vsat_ss=-1000.03                   vsat_ff=-2758.02 vsat_sf=1000.03                    vsat_fs=-1000.03                   wvsat_ss=-2.6e-09 wvsat_ff=0.00508522                 wvsat_sf=2.6e-09                    wvsat_fs=-2.6e-09 lvsat_ss=-4.9e-10                   lvsat_ff=0.000237901                lvsat_sf=4.9e-10 lvsat_fs=-4.9e-10                   pvsat_ss=6.3e-16                    pvsat_ff=-2.5426e-10 pvsat_sf=-6.3e-16                   pvsat_fs=6.3e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.21 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.46085293 lvth0=-3.5855836e-009            wvth0=-2.5374756e-008            pvth0=7.137911e-016 k2=0.021115545                lk2=-2.5584207e-009            wk2=-7.4074707e-009 pk2=1.9505145e-016             minv=-0.79025732                cit=0.0047071352 wcit=-2.695806e-009             voff=-0.19355568                lvoff=-2.3316531e-009 wvoff=6.2710328e-009             pvoff=-1.1883561e-016            eta0=-0.072214321 weta0=1.9057153e-008             etab=-0.043575098               wetab=-3.5788551e-009 u0=0.015174165                wu0=-7.9502993e-011            ua=-2.3207785e-009 lua=4.1059874e-017             wua=1.063767e-017              pua=1.6133951e-024 ub=1.6905843e-018             wub=1.0912485e-025             uc=9.2908642e-011 luc=-1.8011654e-018            wuc=-5.6309452e-017            puc=1.301815e-024 vsat=138833.79                  wvsat=0.00063338744              a0=-3.7689357 la0=-1.9939406e-007            wa0=1.9147626e-006             pa0=-6.1272404e-014 ags=2.7629289                  lags=1.0612622e-008             wags=5.9552827e-008 pags=-2.9290837e-015            keta=-0.53237037                lketa=1.030163e-008 wketa=8.7440889e-008             pketa=-2.4409031e-015            pclm=1.6057928 lpclm=-2.0352482e-008            wpclm=-9.7789759e-007            ppclm=3.9508446e-014 pdiblc2=0.0039674074               lpdiblc2=-8.941037e-011             wpdiblc2=-8.5580444e-010 ppdiblc2=4.8818062e-017             aigbacc=0.015076188                waigbacc=-7.1689126e-011 aigc=0.010503481                laigc=3.3866692e-012             waigc=9.7657768e-012 paigc=-1.7620066e-019            aigsd=0.0099468982               laigsd=-1.1495668e-011 waigsd=-7.0666011e-011            paigsd=3.2079667e-018             bigsd=0.00086753404 wbigsd=-1.0078349e-010            tvoff=-0.000899219               ltvoff=8.6644e-011 wtvoff=1.5106e-009                ptvoff=-5.53421e-017              kt1=-0.30770897 lkt1=2.5841111e-009             wkt1=8.8767065e-008             pkt1=-3.1249354e-015 kt2=-0.087983506               wkt2=4.349409e-009              ua1=1.1554355e-009 lua1=-3.4282991e-017            wua1=-5.2387752e-017            pua1=-1.6355771e-024 ub1=-6.4067874e-019            wub1=-2.5134803e-025            uc1=2.2105679e-010 luc1=-5.8051951e-018            wuc1=2.9270993e-017             puc1=-6.509075e-025 at=129443.41                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.4673854e-010 pcit=8.1914137e-017             lu0=9.4117373e-011             pu0=8.7058878e-018 lub=-2.4490171e-026            pub=-7.0897674e-033            laigbacc=-1.2323729e-010 paigbacc=8.7058878e-018             lbigsd=-1.4898995e-011            pbigsd=4.124872e-018 lkt2=8.6258331e-010             pkt2=-1.2489288e-016            lub1=8.7807268e-027 pub1=1.3965709e-032             lat=-0.0015873796              lvsat=0.00084062967 pvsat=-6.8659594e-011            wat=-0.034682028               pat=1.1818321e-009 letab=7.8076572e-010             petab=8.4122935e-017             leta0=3.0610094e-009 peta0=-7.2413459e-016            lminv=1.499482e-008              wminv=-6.2034136e-008 pminv=2.5433996e-015             vth0_ss=-0.0108247                 vth0_ff=0.0107852 lvth0_ss=4.43812e-10                lvth0_ff=-4.42193e-10               wvth0_ss=3.96894e-09 wvth0_ff=-2.97671e-09               pvth0_ss=-1.62727e-16               pvth0_ff=1.22045e-16 voff_ss=0.0143802                  voff_ff=-0.0106667                 voff_mcl=-0.0109037 voff_mc=0.00835951                 lvoff_ss=-5.8959e-10                lvoff_ff=4.37333e-10 lvoff_mcl=4.47052e-10                lvoff_mc=-3.4274e-10                wvoff_ss=-3.96895e-09 wvoff_ff=-2.2e-15                   wvoff_mcl=5.95342e-09                wvoff_mc=-4.56429e-09 pvoff_ss=1.62727e-16                pvoff_ff=3.1e-22                    pvoff_mcl=-2.4409e-16 pvoff_mc=1.87136e-16                u0_ss=0.000711106                u0_ff=0.000533335 u0_sf=0.000719012                wu0_ss=-1.9e-16                   wu0_ff=1.1e-16 wu0_sf=-1.98447e-10               vsat_ss=-1000.01                   vsat_ff=12091.4 vsat_sf=11666.7                    vsat_fs=-4555.56                   vsat_mc=16703.2 wvsat_ss=2.6e-09                    wvsat_ff=-0.00508522                wvsat_sf=-1.9e-09 wvsat_fs=2.6e-09                    wvsat_mc=-0.00426662                lu0_ss=-2.91555e-11 lu0_ff=-2.18667e-11               lu0_sf=-2.94795e-11               pu0_ss=1.3e-23 pu0_ff=-1.6e-23                   pu0_sf=8.13634e-18                lvsat_ss=-2.8e-10 lvsat_ff=-0.000370923               lvsat_sf=-0.000437333               lvsat_fs=0.000145778 lvsat_mc=-0.000684832               pvsat_ss=-6.3e-17                   pvsat_ff=1.62727e-10 pvsat_sf=1.3e-16                    pvsat_fs=3.7e-17                    pvsat_mc=1.74931e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_mac.22 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.33331005 lvth0=3.8562483e-009             wvth0=-6.0554909e-009            pvth0=-1.0639949e-015 k2=-0.032425692               lk2=-1.1005619e-012            wk2=-2.0217712e-011 pk2=1.6733583e-019             minv=-0.42453                   cit=0.001462963 wcit=-1.5537778e-010            voff=-0.14438889                lvoff=-2.8883421e-008 wvoff=2.647909e-009              pvoff=2.2181564e-017             eta0=0.0072518518 weta0=-6.2151111e-010            etab=-0.055975704               wetab=9.0740622e-010 u0=0.020056926                wu0=-5.9043556e-011            ua=-1.5360414e-009 lua=-5.0886439e-017            wua=1.8604282e-019             pua=-6.9662072e-024 ub=2.0504222e-018             wub=9.3226667e-028             uc=1.2482833e-010 luc=-3.9104259e-017            wuc=9.9259545e-019             puc=-1.9327307e-025 vsat=110740.74                  wvsat=0.0031075556               a0=2.8673811 la0=-7.141216e-007             wa0=9.0352866e-008             pa0=-9.8358479e-014 ags=1.1535045                  lags=7.1999947e-007             wags=1.165353e-008 pags=1.2538332e-014             keta=0.016950323                lketa=-3.5870289e-008 wketa=2.7465313e-009             pketa=-7.2355641e-015            pclm=0.37962963 lpclm=0                          wpclm=1.9422222e-008             ppclm=0 pdiblc2=0.00037156104              lpdiblc2=1.1554369e-009             wpdiblc2=-2.2558551e-011 ppdiblc2=2.0293673e-016             aigbacc=0.012957                   aigc=0.010947941 laigc=-3.6178497e-011            waigc=6.6169369e-012             paigc=3.5102256e-019 aigsd=0.0094977058               laigsd=1.2829566e-010             waigsd=3.9039724e-011 paigsd=-2.0116325e-017            bigsd=0.00036648444              wbigsd=1.5656253e-011 tvoff=0.00231756                 ltvoff=-2.82687e-010              wtvoff=-4.2403e-011 ptvoff=6.85293e-017               kt1=-0.15736741                lkt1=-3.3148323e-012 wkt1=-1.2703068e-009            pkt1=8.4073788e-019             kt2=-0.06021 ua1=1.4600604e-009             lua1=-9.0502337e-017            wua1=2.8927643e-017 pua1=-5.1447263e-024            ub1=-1.1144111e-018            wub1=-6.0247733e-026 uc1=1.0256911e-010             luc1=1.2872267e-017             wuc1=3.9492504e-019 puc1=-3.5527457e-024            at=130000                     jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=0 pcit=0                          lu0=0                          pu0=0 lat=0                          lvsat=0                          pvsat=0 wat=0                          pat=0                          leta0=0 peta0=0                          ags_ff=0.183024                   lags_ff=-1.63989e-07 wags_ff=1.0784e-08                 pags_ff=-9.66244e-15 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_mac.23 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.32168983 lvth0=1.4267971e-008             wvth0=-5.7497722e-009            pvth0=-1.3379189e-015 k2=-0.034041354               lk2=1.4465318e-009             wk2=2.0636638e-010 pk2=-2.0285201e-016            minv=-0.42453                   cit=8.6419753e-005 wcit=-2.1312652e-010            voff=-0.15204641                lvoff=-2.2022286e-008 wvoff=1.1782271e-009             pvoff=1.3390165e-015             eta0=0.0072518518 weta0=-6.2151111e-010            etab=-0.055975704               wetab=9.0740622e-010 u0=0.021237743                wu0=-4.0245607e-010            ua=-1.5629444e-009 lua=-2.6781306e-017            wua=4.5073054e-018             pua=-1.0838059e-023 ub=2.2676811e-018             wub=-2.5439658e-026            uc=7.1641152e-011 luc=8.5514535e-018             wuc=2.3168553e-018             puc=-1.3798099e-024 vsat=110740.74                  wvsat=0.0031075556               a0=2.4025761 la0=-2.9765636e-007            wa0=-2.9047012e-008            pa0=8.623812e-015 ags=1.1513961                  lags=7.2188858e-007             wags=5.492836e-008 pags=-2.6235916e-014            keta=-0.0033042808              lketa=-1.7722164e-008 wketa=-4.1746703e-009            pketa=-1.0341675e-015            pclm=0.29446749 lpclm=7.6305277e-008             wpclm=1.5572306e-008             ppclm=3.4495248e-015 pdiblc2=0.00018729218              lpdiblc2=1.3205418e-009             wpdiblc2=3.0980602e-010 ppdiblc2=-9.4861932e-017            aigbacc=0.012481303                waigbacc=9.6825389e-011 aigc=0.010964676                laigc=-5.1172121e-011            waigc=1.705001e-012 paigc=4.7521171e-018             aigsd=0.009666939                laigsd=-2.3337315e-011 waigsd=7.938917e-012              paigsd=7.7499973e-018             bigsd=0.00027575764 wbigsd=2.6973403e-011             tvoff=0.00231163                 ltvoff=-2.77373e-010 wtvoff=2.61342e-011               ptvoff=7.11996e-018               kt1=-0.13968888 lkt1=-1.5843275e-008            wkt1=-1.4490999e-009            pkt1=1.6103934e-016 kt2=-0.060381058               wkt2=5.4014322e-010             ua1=1.5033473e-009 lua1=-1.2928742e-016            wua1=4.9582026e-017             pua1=-2.3651053e-023 ub1=-1.0770756e-018            wub1=-1.1224085e-025            uc1=1.6079509e-010 luc1=-3.9298205e-017            wuc1=-1.0647109e-017            puc1=6.3409165e-024 at=139911.11                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.2333827e-009 pcit=5.1742872e-017             lu0=-1.0580121e-009            pu0=3.0769761e-016 lub=-1.9466397e-025            pub=2.3629245e-032             laigbacc=4.2622418e-010 paigbacc=-8.6755548e-017            lbigsd=8.1291221e-011             pbigsd=-1.0140166e-017 lkt2=1.5326836e-010             pkt2=-4.8396833e-016            lub1=-3.3452628e-026 pub1=4.6585832e-032             lat=-0.0088803556              lvsat=0 pvsat=0                          wat=0                          pat=0 leta0=0                          peta0=0                          ags_ss=-0.135085 ags_ff=0.202627                   ags_sf=-0.084428                  ags_fs=0.101314 lags_ss=1.21036e-07                lags_ff=-1.81554e-07               lags_sf=7.56475e-08 lags_fs=-9.0777e-08                wags_ss=1.53997e-08                wags_ff=-2.30995e-08 wags_sf=9.62479e-09                wags_fs=-1.15497e-08               pags_ss=-1.37981e-14 pags_ff=2.06971e-14                pags_sf=-8.62381e-15               pags_fs=1.03486e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_mac.24 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.3654446 lvth0=-5.2466585e-009            wvth0=-1.054876e-008             pvth0=8.0242969e-016 k2=-0.030011559               lk2=-3.507566e-010             wk2=-1.8216676e-010 pk2=-2.9566232e-017            minv=-0.42453                   cit=0.0034893954 wcit=-2.7307312e-010            voff=-0.19889571                lvoff=-1.1274963e-009 wvoff=5.5731346e-009             pvoff=-6.2111222e-016            eta0=0.0072518518 weta0=-6.2151111e-010            etab=-0.055975704               wetab=9.0740622e-010 u0=0.018808811                wu0=1.8257553e-010             ua=-1.617289e-009 lua=-2.5436354e-018            wua=-1.9690456e-017            pua=-4.5856883e-026 ub=1.9964359e-018             wub=3.2925149e-026             uc=1.1554479e-010 luc=-1.102957e-017             wuc=-6.0092688e-019            puc=-7.8479058e-026 vsat=110740.74                  wvsat=0.0031075556               a0=1.9918803 la0=-1.1448604e-007            wa0=6.9471795e-008             pa0=-3.5315576e-014 ags=2.6253409                  lags=6.4509211e-008             wags=-2.5022985e-008 pags=9.422384e-015              keta=-0.059812435               lketa=7.480473e-009 wketa=-2.0137906e-009            pketa=-1.9979199e-015            pclm=-0.3541912 lpclm=3.6560705e-007             wpclm=6.201831e-008              ppclm=-1.7265393e-014 pdiblc2=0.0029937954               lpdiblc2=6.8841307e-011             wpdiblc2=1.1470733e-010 ppdiblc2=-7.8479136e-018            aigbacc=0.014090244                waigbacc=-1.2021692e-010 aigc=0.010838498                laigc=5.1031292e-012             waigc=1.7645924e-011 paigc=-2.3575344e-018            aigsd=0.009584091                laigsd=1.3612919e-011 waigsd=4.1258596e-011             paigsd=-7.1105794e-018            bigsd=0.00049846213 wbigsd=6.8819219e-012             tvoff=0.00164385                 ltvoff=2.04541e-011 wtvoff=7.67293e-011               ptvoff=-1.54454e-017              kt1=-0.17556065 lkt1=1.5553181e-010             wkt1=1.0838017e-009             pkt1=-9.6863476e-016 kt2=-0.057542398               wkt2=-6.1619905e-011            ua1=1.6650489e-009 lua1=-2.0140633e-016            wua1=-3.7594673e-017            pua1=1.5229755e-023 ub1=-1.6172312e-018            wub1=3.3640185e-026             uc1=4.4309416e-011 luc1=1.2654404e-017             wuc1=6.8047266e-018             puc1=-1.442602e-024 at=178199.88                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=-2.8434441e-010 pcit=7.8479058e-017             lu0=2.5291687e-011             pu0=4.6773518e-017 lub=-7.3688603e-026            pub=-2.4014592e-033            laigbacc=-2.9136323e-010 paigbacc=1.0045319e-017             lbigsd=-1.8034981e-011            pbigsd=-1.1793654e-018 lkt2=-1.1127744e-009            pkt2=-2.1558197e-016            lub1=2.0745679e-025 pub1=-1.8477109e-032            lat=-0.025957145               lvsat=0 pvsat=0                          wat=-0.0032846802              pat=1.4649674e-009 leta0=0                          peta0=0                          ags_ss=0.167166 ags_ff=-0.266186                  ags_sf=0.116056                   ags_fs=-0.133093 lags_ss=-1.37682e-08               lags_ff=2.75365e-08                lags_sf=-1.37682e-08 lags_fs=1.37683e-08                wags_ss=-1.9057e-08                wags_ff=3.03451e-08 wags_sf=-1.32303e-08               wags_fs=1.51726e-08                pags_ss=1.56958e-15 pags_ff=-3.13917e-15               pags_sf=1.56958e-15                pags_fs=-1.56958e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_mac.25 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.33796819 lvth0=5.783411e-010              wvth0=-5.5008645e-009            pvth0=-2.6772417e-016 k2=-0.028414861               lk2=-6.8925657e-010            wk2=-5.4796804e-010 pk2=4.7983639e-017             minv=-0.42453                   cit=0.00095859271 wcit=1.5749418e-010             voff=-0.19093415                lvoff=-2.8153472e-009 wvoff=2.4314554e-009             pvoff=4.4923765e-017             eta0=0.0072518518 weta0=-6.2151111e-010            etab=-0.055976141               wetab=9.0748921e-010 u0=0.019380812                wu0=4.1182202e-010             ua=-1.6422933e-009 lua=2.7572903e-018             wua=-3.4197675e-017            pua=3.0296735e-024 ub=1.7603448e-018             wub=4.2516169e-026             uc=9.8822252e-011 luc=-7.4843914e-018            wuc=-1.2958938e-018            puc=6.8853936e-026 vsat=114750.16                  wvsat=0.0010164811               a0=4.9722399 la0=-7.4632226e-007            wa0=-3.754963e-007             pa0=5.9017659e-014 ags=2.9432071                  lags=-2.8784266e-009            wags=1.9687351e-008 pags=-5.6207295e-017            keta=0.035075365                lketa=-1.2635741e-008 wketa=-1.3942214e-008            pketa=5.30906e-016               pclm=1.4866549 lpclm=-2.4652322e-008            wpclm=-3.267866e-008             ppclm=2.8103647e-015 pdiblc2=0.0035359202               lpdiblc2=-4.6089134e-011            wpdiblc2=1.3071461e-010 ppdiblc2=-1.1241456e-017            aigbacc=0.012446008                waigbacc=-2.2458871e-011 aigc=0.01094271                 laigc=-1.6989934e-011            waigc=2.1574556e-012 paigc=9.260208e-019              aigsd=0.0096965317               laigsd=-1.0224521e-011 waigsd=9.3680338e-012             paigsd=-3.4978024e-019            bigsd=0.00038847748 wbigsd=1.5509395e-012             tvoff=0.00170806                 ltvoff=6.84197e-012 wtvoff=1.3909e-011                ptvoff=-2.12753e-018              kt1=-0.16577471 lkt1=-1.9190864e-009            wkt1=-3.5326268e-009            pkt1=1.0048094e-017 kt2=-0.053410811               wkt2=-3.0848778e-009            ua1=1.0858386e-009 lua1=-7.8613748e-017            wua1=3.1724474e-017             pua1=5.3409591e-025 ub1=-9.1299643e-019            wub1=-5.3423196e-026            uc1=8.8630217e-011 luc1=3.2583939e-018             wuc1=4.24206e-018               puc1=-8.9931671e-025 at=53013.222                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=2.5218575e-010 pcit=-1.2801211e-017            lu0=-9.5972562e-011            pu0=-1.8267371e-018 lub=-2.363729e-026             pub=-4.4347555e-033            laigbacc=5.7214824e-011 paigbacc=-1.0679386e-017            lbigsd=5.2817635e-012             pbigsd=-4.9197121e-020 lkt2=-1.9886707e-009            pkt2=4.253487e-016              lub1=5.8159008e-026 pub1=-1.9672553e-035            lat=0.00058242554              lvsat=-0.00084999803 pvsat=4.4330778e-010             wat=0.0035800407               pat=9.6465404e-012 letab=9.2682013e-014             petab=-1.7592883e-020            leta0=0 peta0=0                          ua_ss=3.36214e-11                lua_ss=-7.12774e-18 wua_ss=-9.27951e-18               pua_ss=1.96726e-24                vsat_ss=4651.38 vsat_ff=-5814.23                   vsat_sf=2325.69                    vsat_fs=-2907.11 wvsat_ss=-0.000530258               wvsat_ff=0.000662822                wvsat_sf=-0.000265129 wvsat_fs=0.000331411                ags_ss=0.171993                   ags_ff=-0.229324 ags_sf=0.0859965                  ags_fs=-0.114662                  lags_ss=-1.47914e-08 lags_ff=1.97219e-08                lags_sf=-7.3957e-09                lags_fs=9.86093e-09 wags_ss=-1.96072e-08               wags_ff=2.61429e-08                wags_sf=-9.8036e-09 wags_fs=1.30715e-08                pags_ss=1.68622e-15                pags_ff=-2.24829e-15 pags_sf=8.43109e-16                pags_fs=-1.12415e-15               lvsat_ss=-0.000986093 lvsat_ff=0.00123262                 lvsat_sf=-0.000493046               lvsat_fs=0.000616308 pvsat_ss=1.12415e-10                pvsat_ff=-1.40518e-10               pvsat_sf=5.62073e-11 pvsat_fs=-7.02591e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_mac.26 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.3301285 lvth0=1.2525545e-009             wvth0=-1.1317632e-008            pvth0=2.3251789e-016 k2=-0.02451211                lk2=-1.0248932e-009            wk2=8.7524126e-011 pk2=-6.6686869e-018            minv=-0.42453                   cit=0.0023352547 wcit=1.0157283e-010             voff=-0.20588095                lvoff=-1.5299224e-009 wvoff=3.69158e-009               pvoff=-6.3446953e-017            eta0=0.009618107 weta0=-8.912642e-010             etab=-0.087079114               wetab=2.8958135e-009 u0=0.017843298                wu0=7.1967965e-010             ua=-1.9732314e-009 lua=3.1217962e-017             wua=-1.3845836e-017            pua=1.2794154e-024 ub=1.7635317e-018             wub=3.2162121e-026             uc=2.3031584e-011 luc=-9.6639403e-019            wuc=6.3699494e-018             puc=-5.9040858e-025 vsat=99488.669                  wvsat=0.0035691502               a0=6.8264815 la0=-9.0578704e-007            wa0=-4.7098889e-007            pa0=6.7230022e-014 ags=2.909737                   lags=0                          wags=1.9033778e-008 pags=0                          keta=0.015374486                lketa=-1.0941465e-008 wketa=-2.3716691e-008            pketa=1.371511e-015              pclm=1.4484568 lpclm=-2.1367284e-008            wpclm=8.0925926e-009             ppclm=-6.9596296e-016 pdiblc2=0.0035967078               lpdiblc2=-5.1316872e-011            wpdiblc2=2.6975309e-011 ppdiblc2=-2.3198765e-018            aigbacc=0.016196533                waigbacc=-6.1789642e-010 aigc=0.010853664                laigc=-9.3319237e-012            waigc=2.71609e-011 paigc=-1.2242754e-018            aigsd=0.0096446803               laigsd=-5.7652959e-012 waigsd=-1.3516423e-011            paigsd=1.618283e-018              bigsd=0.00047987472 wbigsd=-9.6178316e-012            tvoff=0.00183695                 ltvoff=-4.2426e-012 wtvoff=-6.45682e-012              ptvoff=-3.76067e-019              kt1=-0.19030513 lkt1=1.9052993e-010             wkt1=-2.8015244e-009            pkt1=-5.2826721e-017 kt2=-0.091507626               wkt2=3.468496e-009              ua1=1.1033926e-009 lua1=-8.0123392e-017            wua1=-4.9334596e-017            pua1=7.5051759e-024 ub1=-1.4972618e-018            wub1=9.680014e-026              uc1=1.2938272e-011 luc1=9.7679012e-018             wuc1=6.733037e-018              puc1=-1.1135407e-024 at=74787.869                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.3379282e-010 pcit=-7.9919747e-018            lu0=3.6253601e-011             pu0=-2.8302494e-017 lub=-2.3911362e-026            pub=-3.5443074e-033            laigbacc=-2.6533035e-010 paigbacc=4.0528243e-017             lbigsd=-2.5783994e-012            pbigsd=9.113172e-019 lkt2=1.2876554e-009             pkt2=-1.3824144e-016            lub1=1.0840583e-025 pub1=-1.2938879e-032            lat=-0.0012901941              lvsat=0.00046249065 pvsat=2.2377824e-010             wat=0.00055430892              pat=2.6985947e-010 letab=2.6749484e-009             petab=-1.7101348e-016            leta0=-2.0349794e-010 peta0=2.3198765e-017             ua_ss=-6.88066e-11               lua_ss=1.68107e-18 wua_ss=1.89906e-17                pua_ss=-4.63974e-25               vsat_ss=-13913.5 vsat_ff=15617.3                    vsat_sf=-10506.2                   vsat_fs=12541.2 wvsat_ss=0.00158615                 wvsat_ff=-0.00178037                wvsat_sf=0.0011977 wvsat_fs=-0.00142969                lvsat_ss=0.000610494                lvsat_ff=-0.000610494 lvsat_sf=0.000610494                lvsat_fs=-0.000712243               pvsat_ss=-6.95963e-11 pvsat_ff=6.95965e-11                pvsat_sf=-6.95963e-11               pvsat_fs=8.11957e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_mac.27 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.29189446 lvth0=3.1642562e-009             wvth0=-6.1964594e-009            pvth0=-2.354077e-017 k2=-0.024479344               lk2=-1.0265315e-009            wk2=1.4680021e-009 pk2=-7.5692587e-017            minv=-0.42453                   cit=0.0023882922 wcit=-5.3826531e-010            voff=-0.19220818                lvoff=-2.2135607e-009 wvoff=3.4107914e-009             pvoff=-4.9407521e-017            eta0=-0.0184107 weta0=1.7846864e-009             etab=-0.050418063               wetab=-2.6861957e-009 u0=0.022913189                wu0=4.3056909e-010             ua=-2.4743563e-009 lua=5.6274206e-017             wua=1.1098369e-016             pua=-4.962061e-024 ub=2.9608744e-018             wub=-1.4550313e-025            uc=1.1303704e-010 luc=-5.4666667e-018            wuc=-5.4382222e-018            puc=4.8567097e-039 vsat=-10215.723                 wvsat=0.018648492                a0=-30.942406 la0=9.8265732e-007             wa0=5.0221009e-006             pa0=-2.0742447e-013 ags=2.909737                   lags=0                          wags=1.9033778e-008 pags=0                          keta=-0.40647737                lketa=1.0151128e-008 wketa=4.717442e-008              pketa=-2.1730445e-015            pclm=0.83003353 lpclm=9.553879e-009              wpclm=-2.5590489e-008            ppclm=9.8819112e-016 pdiblc2=0.00029259259              lpdiblc2=1.1388889e-010             wpdiblc2=-1.9422222e-011 ppdiblc2=1.0864276e-031             aigbacc=0.00036642387              waigbacc=1.8498803e-009 aigc=0.011086204                laigc=-2.0958938e-011            waigc=-2.3968824e-011 paigc=1.3322108e-018             aigsd=0.0087006767               laigsd=4.143488e-011 waigsd=1.2648786e-010             paigsd=-5.381931e-018             bigsd=8.6761222e-005 wbigsd=4.7544701e-011             tvoff=0.000568066                ltvoff=5.92016e-011 wtvoff=1.93147e-010               ptvoff=-1.03563e-017              kt1=-0.25867398 lkt1=3.6089722e-009             wkt1=1.4480484e-008             pkt1=-9.1692712e-016 kt2=-0.07538935                wkt2=2.1281792e-009             ua1=-9.1726746e-010 lua1=2.0909611e-017             wua1=6.6708059e-017             pua1=1.7030432e-024 ub1=1.6415121e-018             wub1=-1.9473238e-025            uc1=3.6892181e-010 luc1=-8.0312757e-018            wuc1=-2.969442e-017             puc1=7.078321e-025 at=48012.229                  jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=1.3114095e-010 pcit=2.3999932e-017             lu0=-2.1724095e-010            pu0=-1.3846965e-017 lub=-8.3778498e-026            pub=5.3389554e-033             laigbacc=5.261751e-010 paigbacc=-8.2860595e-017            lbigsd=1.7077276e-011             pbigsd=-1.9468094e-018 lkt2=4.8174156e-010             pkt2=-7.1225605e-017            lub1=-4.8532864e-026 pub1=1.6377465e-033             lat=4.8587885e-005             lvsat=0.0059477103 pvsat=-5.3018885e-010            wat=0.0075286283               pat=-7.88565e-011 letab=8.418958e-010              petab=1.0808698e-016             leta0=1.1979424e-009 peta0=-1.1059876e-016            u0_sf=-0.000320576               wu0_sf=8.8479e-11 ua_ss=-3.51853e-11               lua_ss=3.3e-24                    wua_ss=9.71112e-18 pua_ss=4.7e-30                    vsat_ss=-1703.7                    vsat_ff=26691.3 vsat_sf=1703.7                     vsat_fs=-1703.7                    wvsat_ss=0.00019422 wvsat_ff=-0.00304281                wvsat_sf=-0.00019422                wvsat_fs=0.00019422 ua1_sf=-9.61728e-11               lua1_sf=4.80864e-18                wua1_sf=2.65437e-17 pua1_sf=-1.32719e-24               at_ss=32057.6                    lu0_sf=1.60288e-11 pu0_sf=-4.42395e-18               lat_ss=-0.00160288                lvsat_ss=1.6e-10 lvsat_ff=-0.0011642                 lvsat_sf=-1.6e-10                   lvsat_fs=1.6e-10 pvsat_ss=6e-18                      pvsat_ff=1.32719e-10                pvsat_sf=-6e-18 pvsat_fs=6e-18                      wat_ss=-0.0088479                 pat_ss=4.42395e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_mac.28 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.4934563 lvth0=-5.0997792e-009            wvth0=-3.4373285e-008            pvth0=1.1317091e-015 k2=-0.019937418               lk2=-1.2127504e-009            wk2=3.9231474e-009 pk2=-1.7635354e-016            minv=-1.2440694                 cit=-0.0034607202 wcit=-4.414779e-010             voff=-0.23475283                lvoff=-4.6923007e-010 wvoff=1.7641446e-008             pvoff=-6.3286435e-016            eta0=0.005144856 weta0=-2.2939803e-009            etab=-0.053893472               wetab=-7.3098416e-010 u0=0.020742333                wu0=-1.6163173e-009            ua=-2.5235332e-009 lua=5.829046e-017              wua=6.6597978e-017             pua=-3.1422467e-024 ub=2.7043992e-018             wub=-1.7068805e-025            uc=-7.1390947e-011 luc=2.0948807e-018             wuc=-1.0962765e-017            puc=2.2650627e-025 vsat=147787.12                  wvsat=-0.0018377314              a0=3.7798542 la0=-4.4095533e-007            wa0=-1.6870337e-007            pa0=5.398508e-015 ags=2.7178292                  lags=7.8682206e-009             wags=7.2000336e-008 pags=-2.1716289e-015            keta=-0.044320988               lketa=-4.697284e-009 wketa=-4.7260741e-008            pketa=1.698797e-015              pclm=-2.1629553 lpclm=1.3226642e-007             wpclm=6.2276909e-008             ppclm=-2.6143722e-015 pdiblc2=0.0011872428               lpdiblc2=7.720823e-011              wpdiblc2=-8.8479012e-011 ppdiblc2=2.8313284e-018             aigbacc=0.016382185                waigbacc=-4.3214444e-010 aigc=0.010047488                laigc=2.162841e-011              waigc=1.3561976e-010 paigc=-5.2109212e-018            aigsd=0.010016824                laigsd=-1.2527166e-011 waigsd=-8.9965586e-011            paigsd=3.4926602e-018             bigsd=0.00050136063 wbigsd=2.8036787e-013             tvoff=0.0069069                  ltvoff=-2.00691e-010 wtvoff=-6.4389e-010               ptvoff=2.39623e-017               kt1=0.19196238 lkt1=-1.4867119e-008            wkt1=-4.9142227e-008            pkt1=1.691604e-015 kt2=-0.080679621               wkt2=2.3335368e-009             ua1=6.7513086e-010 lua1=-4.437872e-017             wua1=8.0176331e-017             pua1=1.150844e-024 ub1=-1.2591072e-018            wub1=-8.0661784e-026            uc1=5.0225514e-010 luc1=-1.3497942e-017            wuc1=-4.8339753e-017            puc1=1.4722908e-024 at=-50946.511                 jtsswgs='4.52e-005*(1+1.57*iboffn_flag)' jtsswgd='4.52e-005*(1+1.57*iboffn_flag)'                                   lcit=3.7095045e-010 pcit=2.0031648e-017             lu0=-1.2823585e-010            pu0=7.0075378e-017 lub=-7.3263014e-026            pub=6.3715371e-033             laigbacc=-1.3047111e-010 paigbacc=1.0702421e-017             lbigsd=7.8699753e-014             pbigsd=-8.9717718e-021 lkt2=6.986427e-010              pkt2=-7.9645268e-017            lub1=7.0392525e-026 pub1=-3.0391479e-033            lat=0.0041058963               lvsat=-0.0005304062 pvsat=3.0974631e-010             wat=0.015105591                pat=-3.8951198e-010 letab=9.8438756e-010             petab=2.7923305e-017             leta0=2.3216461e-010 peta0=5.6626568e-017             lminv=3.3601116e-008             wminv=6.3217998e-008 pminv=-2.5919379e-015            vth0_ss=0.00605761                 lvth0_ss=-2.48362e-10 wvth0_ss=-6.90568e-10               pvth0_ss=2.83133e-17                voff_ff=-0.0181728 voff_mcl=0.0181728                  voff_mc='-0.0139325+0.00500412'    lvoff_ff=7.45086e-10 lvoff_mcl=-7.45086e-10               lvoff_mc='5.71233e-10-2.05169e-10'  wvoff_ff=2.0717e-09 wvoff_mcl=-2.0717e-09                wvoff_mc='1.58831e-09-1.38114e-09'  pvoff_ff=-8.49399e-17 pvoff_mcl=8.49399e-17                pvoff_mc='-6.51206e-17+5.66266e-17' u0_ss=0.00121152 u0_ff=0.000908642                u0_sf=0.000320576                wu0_ss=-1.38114e-10 wu0_ff=-1.03585e-10               wu0_sf=-8.8479e-11                ua_ss=-1.60288e-10 lua_ss=5.12922e-18                wua_ss=4.42395e-17                pua_ss=-1.41566e-24 vsat_ss=-1703.71                   vsat_ff=-10790.1                   vsat_sf=19876.5 vsat_fs=-7761.32                   vsat_mc=-10390.1                   wvsat_ss=0.000194222 wvsat_ff=0.00123007                 wvsat_sf=-0.00226593                wvsat_fs=0.00088479 wvsat_mc=0.00321114                 ua1_sf=9.61728e-11                lua1_sf=-3.07753e-18 wua1_sf=-2.65437e-17               pua1_sf=8.49399e-25                at_ss=68024.7 at_sf=15012.3                    lu0_ss=-4.96724e-11               lu0_ff=-3.72543e-11 lu0_sf=-1.02584e-11               pu0_ss=5.66266e-18                pu0_ff=4.24699e-18 pu0_sf=2.83133e-18                lat_ss=-0.00307753                lat_sf=-0.000615506 lvsat_ss=1.4e-10                    lvsat_ff=0.000372543                lvsat_sf=-0.000745086 lvsat_fs=0.000248362                lvsat_mc=0.000425995                pvsat_ss=1.6e-17 pvsat_ff=-4.24699e-11               pvsat_sf=8.49399e-11                pvsat_fs=-2.83133e-11 pvsat_mc=-1.31657e-10               wat_ss=-0.0187748                 wat_sf=-0.00414341 pat_ss=8.49398e-10                pat_sf=1.6988e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model pch_mac.global pmos ( modelid=2                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag'                 permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=2.18e-009                  toxm=2.18e-009                  dtox=6.63e-010 epsrox=3.9                        wint=0                          lint=0 ll=0                          wl=0                          lln=1 wln=1                          lw=0                          ww=0 lwn=1                          wwn=1                          lwl=0 wwl=0                          llc=0                          wlc=0 lwc=0                          wwc=0                          lwlc=0 wwlc=0                          xl=-3e-009                    xw=6e-009 dlc=6.67e-009                  dwc=0                          xpart=1 toxref=3e-009                     dlcig=2.5e-009                   k1=0.35 k3=0                          k3b=1.5                        w0=0 dvt0=1.166                      dvt1=0.9918                     dvt2=2.22e-016 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.2                        minv=-0.33                      voffl=0 dvtp0=1.07e-007                  dvtp1=0.5                        lpe0=1.335e-008 lpeb=4.44089e-021               xj=8.5e-008                   ngate=4.5674e+019 ndep=6e+017                     nsd=1e+020                     phin=0.2 cdsc=0                          cdscb=0                          cdscd=0 nfactor=0.7                        ud=0                          lud=0 wud=0                          pud=0                          a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=2.1 delta=0.018814                   pscbe1=9.264e+008                 pscbe2=1e-020 fprout=200                        pdits=0                          pditsd=0 pditsl=0                          rsh=16.7                       rdsw=160 prwg=0                          prwb=0                          wr=1 alpha0=1.8425e-006                alpha1=2                          beta0=19 agidl=6.03e-007                  bgidl=2.68e+009                  cgidl=0.2 egidl=0.001                      bigbacc=0.006993                   cigbacc=0.245 nigbacc=7.236                      aigbinv=0.008351                   bigbinv=0.001095 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1.697 bigc=0.001431                   cigc=0.15259                    cigsd=0.0011 nigc=0.9942                     poxedge=1                          pigcd=3.332 ntox=1                          xrcrg1=12                         xrcrg2=1 vfbsdoff=0.01                       lvfbsdoff=0                          wvfbsdoff=0 pvfbsdoff=0                          cgso=5.02e-011                  cgdo=5.02e-011 cgbo=0                          cgdl=6.0796e-011                cgsl=6.0796e-011 clc=0                          cle=0.6                        cf='9e-011+0.92e-10*ccoflag' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=6                          noff=2.289                      voffcv=-0.078645 tvfbsdoff=0.1                        ltvfbsdoff=0                          wtvfbsdoff=0 ptvfbsdoff=0                          kt1l=0                          prt=0 fnoimod=1.000000e+00               tnoimod=1                          em=2.000000e+07 ef=1.040000e+00               noia=0                          noib=0 noic=0                          lintnoi=-4.230000e-08              jss=4.45e-07 jsd=4.45e-07                   jsws=9.12e-14                   jswd=9.12e-14 jswgs=9.12e-14                   jswgd=9.12e-14                   njs=1.02 njd=1.02                       ijthsfwd=0.01                       ijthdfwd=0.01 ijthsrev=0.01                       ijthdrev=0.01                       bvs=7.43 bvd=7.43                       xjbvs=1                          xjbvd=1 njtsswg=8.7214                     xtsswgs=0.1                        xtsswgd=0.1 tnjtsswg=1                          vtsswgs=1.338                      vtsswgd=1.338 pbs=0.789                      pbd=0.789                      cjs=0.001514 cjd=0.001514                   mjs=0.4                        mjd=0.4 pbsws=0.770                      pbswd=0.770                      cjsws=1.129e-010 cjswd=1.129e-010                 mjsws=0.277                      mjswd=0.277 pbswgs=0.941                      pbswgd=0.941                      cjswgs=2.08e-010 cjswgd=2.08e-010                  mjswgs=0.704                      mjswgd=0.704 tpb=0.00105                    tcj=0.00076                    tpbsw=0.00097 tcjsw=0.00034                    tpbswg=0.00202                    tcjswg=0.00157 xtis=3                          xtid=3                          dmcg=3.75e-008 dmci=3.75e-008                  dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=-5.1e-009 rshg=14.4                       gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          lnfactor=0 pnfactor=0                          wnfactor=0                          pk2we=0 lk2we=0                          wk2we=0                          k2we=0.0000 pku0we=4.5e-18                    wku0we=-1.0e-10                   lku0we=-2e-11 ku0we=-0.0007                    pkvth0we=1e-019                     wkvth0we=-1e-011 lkvth0we=10e-012                    kvth0we=-0.0004346                 wec=-7896.1 web=2251.7                     scref=1e-6                       rnoia=0 rnoib=0                          tnoia=0                          wpemod=1 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.2                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.4 bidirectionflag='bidirectionflag_mos' iboffn_flag='iboffn_flag' iboffp_flag='iboffp_flag' sigma_factor='sigma_factor' ccoflag='ccoflag' rcoflag='rcoflag' rgflag='rgflag' mismatchflag='mismatchflag_mos' globalflag='globalflag_mos' totalflag='totalflag_mos' designflag='designflag_mos' global_factor='global_factor' local_factor='local_factor' sigma_factor_flicker='sigma_factor_flicker' noiseflag='noiseflagp' noiseflag_mc='noiseflagp_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w11='2.3875*0.35355' w12='0.70711*0.35355' w13='0.54772*0.32451' w14='0.54772*-0.16328' w15='0.54772*0.12195' w16='0.54772*0.66871' w17='0.54772*0.32929' w18='0.54772*-0.21807' w19='0' w20='0' tox_c='toxp'                     dxl_c='dxlp'                     dxw_c='dxwp' cj_c='cjp'                      cjsw_c='cjswp'                    cjswg_c='cjswgp' cgo_c='cgop'                     cgl_c='cglp'                     ddlc_c='ddlcp' cf_c='cfp'                      ntox_c='ntoxp'                    dvth_c='dvthp' dlvth_c='dlvthp'                   dwvth_c='dwvthp'                   dpvth_c='dpvthp' dk2_c='dk2p'                     dlk2_c='dlk2p'                    dwk2_c='dwk2p' dpk2_c='dpk2p'                    deta0_c='deta0p'                   dleta0_c='dleta0p' dweta0_c='dweta0p'                  dpeta0_c='dpeta0p'                  dvoff_c='dvoffp' dlvoff_c='dlvoffp'                  dwvoff_c='dwvoffp'                  dpvoff_c='dpvoffp' dcit_c='dcitp'                    dlcit_c='dlcitp'                   dwcit_c='dwcitp' dpcit_c='dpcitp'                   dnfactor_c='dnfactorp'                dlnfactor_c='dlnfactorp' dwnfactor_c='dwnfactorp'               dpnfactor_c='dpnfactorp'               du0_c='du0p' dlu0_c='dlu0p'                    dwu0_c='dwu0p'                    dpu0_c='dpu0p' dpclm_c='dpclmp'                   dlpclm_c='dlpclmp'                  dwpclm_c='dwpclmp' dppclm_c='dppclmp'                  dpdiblc2_c='dpdiblc2p'                dlpdiblc2_c='dlpdiblc2p' dvsat_c='dvsatp'                   dlvsat_c='dlvsatp'                  dwvsat_c='dwvsatp' dpvsat_c='dpvsatp'                  da0_c='da0p'                     dags_c='dagsp' dwags_c='dwagsp'                   dlags_c='dlagsp'                   dpags_c='dpagsp' jtsswg_c='jtsswgp'                  dminv_c='dminvp'                   dat_c='datp' dlat_c='dlatp'                    dwat_c='dwatp'                    dpat_c='dpatp' dua1_c='dua1p'                    dlua1_c='dlua1p'                   dwua1_c='dwua1p' dpua1_c='dpua1p'                   dketa_c='dketap'                   dlketa_c='dlketap' dwketa_c='dwketap'                  dpketa_c='dpketap'                  ss_flag_c='ss_flagp' ff_flag_c='ff_flagp'                 sf_flag_c='sf_flagp'                 fs_flag_c='fs_flagp' monte_flag_c='monte_flagp'             c1f_c='c1fp'                     c2f_c='c2fp' c3f_c='c3fp' global_mc='global_mc_flag' tox_g='toxp_ms_global'           dxl_g='dxlp_ms_global'           dxw_g='dxwp_ms_global' cj_g='cjp_ms_global'            cjsw_g='cjswp_ms_global'          cjswg_g='cjswgp_ms_global' cgo_g='cgop_ms_global'           cgl_g='cglp_ms_global'           cf_g='cfp_ms_global' ntox_g='ntoxp_ms_global'          dvth_g='dvthp_ms_global'          dlvth_g='dlvthp_ms_global' dwvth_g='dwvthp_ms_global'         dpvth_g='dpvthp_ms_global'         dk2_g='dk2p_ms_global' dlk2_g='dlk2p_ms_global'          deta0_g='deta0p_ms_global'         dlvoff_g='dlvoffp_ms_global' dpvoff_g='dpvoffp_ms_global'        du0_g='du0p_ms_global'           dlu0_g='dlu0p_ms_global' dwu0_g='dwu0p_ms_global'          dpu0_g='dpu0p_ms_global'          dlpclm_g='dlpclmp_ms_global' dpdiblc2_g='dpdiblc2p_ms_global'      dvsat_g='dvsatp_ms_global'         dlvsat_g='dlvsatp_ms_global' dwvsat_g='dwvsatp_ms_global'        dpvsat_g='dpvsatp_ms_global'        dags_g='dagsp_ms_global' dwags_g='dwagsp_ms_global'         dminv_g='dminvp_ms_global'         dat_g='datp_ms_global' dpat_g='dpatp_ms_global'          dua1_g='dua1p_ms_global'          dpua1_g='dpua1p_ms_global' dketa_g='dketap_ms_global'         dpketa_g='dpketap_ms_global'        ss_flag_g='ss_flagp_ms_global' ff_flag_g='ff_flagp_ms_global'       monte_flag_g='monte_flagp_ms_global' sf_flag_g='sf_flagp_ms_global'       fs_flag_g='fs_flagp_ms_global' weight1=-3.6045455 weight2=2.1424476 weight3=1.2984615 weight4=-0.6993007 weight5=-0.48664336 tox_1=4.007296e-012 tox_2=-1.002299e-011 tox_3=-3.0894969e-012 tox_4=3.7476963e-011 tox_5=7.4492926e-013 dxl_1=9.0730909e-011 dxl_2=-2.2692977e-010 dxl_3=-6.995093e-011 dxl_4=-8.4852915e-010 dxl_5=1.6865983e-011 dxw_1=-6.8642931e-010 dxw_2=-8.2779917e-010 dxw_3=2.4601975e-010 dxw_4=-1.2698987e-025 dxw_5=-5.8968941e-009 cj_1=9.9548e-006 cj_2=-3.0995e-006 cj_3=-4.9466e-006 cj_4=-1.1157e-022 cj_5=-9.4661e-007 cjsw_1=7.4233e-013 cjsw_2=-2.3113e-013 cjsw_3=-3.6887e-013 cjsw_4=-3.344e-028 cjsw_5=-7.059e-014 cjswg_1=1.3676e-012 cjswg_2=-4.2583e-013 cjswg_3=-6.7958e-013 cjswg_4=-6.1607e-028 cjswg_5=-1.3005e-013 cgo_1=-3.3007e-013 cgo_2=1.0277e-013 cgo_3=1.6401e-013 cgo_4=-4.5203e-028 cgo_5=3.1387e-014 cgl_1=-3.9974e-013 cgl_2=1.2446e-013 cgl_3=1.9863e-013 cgl_4=-3.0195e-028 cgl_5=3.8012e-014 cf_1=-5.9176e-013 cf_2=1.8425e-013 cf_3=2.9405e-013 cf_4=-1.0063e-028 cf_5=5.6272e-014 ntox_1=0.018786 ntox_2=-0.0058493 ntox_3=-0.0093349 ntox_4=-8.4625e-018 ntox_5=-0.0017864 dvth_1=-0.0026306 dvth_2=-0.0036774 dvth_3=0.0011994 dvth_4=1.2765e-018 dvth_5=0.00083771 dlvth_1=-1.6816e-010 dlvth_2=-1.8183e-010 dlvth_3=-6.6104e-012 dlvth_4=-6.4945e-026 dlvth_5=4.2968e-011 dwvth_1=-1.5852e-010 dwvth_2=-8.8382e-011 dwvth_3=9.9465e-011 dwvth_4=-1.8203e-025 dwvth_5=3.4862e-011 dpvth_1=-1.9802e-017 dpvth_2=-4.2262e-018 dpvth_3=1.0779e-017 dpvth_4=1.7263e-033 dpvth_5=3.2574e-018 dk2_1=0.00065287 dk2_2=0.0014524 dk2_3=-0.00011719 dk2_4=-2.8764e-020 dk2_5=-0.00027453 dlk2_1=9.7054e-012 dlk2_2=-3.5921e-012 dlk2_3=1.6826e-011 dlk2_4=4.7997e-027 dlk2_5=5.8634e-014 deta0_1=-0.00018786 deta0_2=5.8493e-005 deta0_3=9.3349e-005 deta0_4=8.4625e-020 deta0_5=1.7864e-005 dlvoff_1=-1.5151e-011 dlvoff_2=6.1206e-012 dlvoff_3=-4.5752e-011 dlvoff_4=-9.7959e-028 dlvoff_5=-9.7498e-013 dpvoff_1=-3.7572e-018 dpvoff_2=1.1699e-018 dpvoff_3=1.867e-018 dpvoff_4=1.6925e-033 dpvoff_5=3.5728e-019 du0_1=4.1979e-005 du0_2=0.00011954 du0_3=-1.0175e-005 du0_4=-3.3672e-020 du0_5=-2.1255e-005 dlu0_1=3.6788e-012 dlu0_2=9.9828e-012 dlu0_3=2.1279e-012 dlu0_4=-3.514e-027 dlu0_5=-2.0292e-012 dwu0_1=6.5311e-012 dwu0_2=1.0847e-011 dwu0_3=-1.7907e-012 dwu0_4=1.082e-027 dwu0_5=-2.4387e-012 dpu0_1=-2.8565e-019 dpu0_2=9.1961e-019 dpu0_3=3.6792e-019 dpu0_4=4.8523e-036 dpu0_5=-9.5417e-020 dpu0_max=-3e-018 dlpclm_1=2.1568e-010 dlpclm_2=-7.9824e-011 dlpclm_3=3.7392e-010 dlpclm_4=1.6123e-026 dlpclm_5=1.303e-012 dpdiblc2_1=-1.8786e-005 dpdiblc2_2=5.8493e-006 dpdiblc2_3=9.3349e-006 dpdiblc2_4=-1.8079e-021 dpdiblc2_5=1.7864e-006 dvsat_1=1382.9 dvsat_2=-440.07 dvsat_3=-326.33 dvsat_4=1.3085e-012 dvsat_5=-115.14 dlvsat_1=8.317e-006 dlvsat_2=7.2783e-005 dlvsat_3=4.9545e-006 dlvsat_4=2.0797e-021 dlvsat_5=-1.0582e-005 dwvsat_1=0.00030526 dwvsat_2=-0.0001036 dwvsat_3=0.00017305 dwvsat_4=-6.4883e-019 dwvsat_5=-1.4305e-005 dpvsat_1=2.0496e-012 dpvsat_2=1.9229e-011 dpvsat_3=-7.1398e-013 dpvsat_4=-1.972e-027 dpvsat_5=-3.4999e-012 dags_1=0.056196 dags_2=0.040452 dags_3=-0.020671 dags_4=5.8482e-017 dags_5=-0.01278 dwags_1=-1.3432e-009 dwags_2=-3.644e-009 dwags_3=-1.6269e-009 dwags_4=4.0421e-025 dwags_5=4.6881e-010 dminv_1=-0.01315 dminv_2=0.0040945 dminv_3=0.0065344 dminv_4=-3.8931e-018 dminv_5=0.0012505 dat_1=1570.7 dat_2=-498.56 dat_3=-419.68 dat_4=-1.7221e-013 dat_5=-133 dpat_1=1.6176e-012 dpat_2=-5.9868e-013 dpat_3=2.8044e-012 dpat_4=4.5526e-028 dpat_5=9.7724e-015 dua1_1=2.957e-012 dua1_2=-9.8405e-013 dua1_3=9.3609e-013 dua1_4=-1.9986e-027 dua1_5=-1.7213e-013 dpua1_1=1.348e-026 dpua1_2=-4.989e-027 dpua1_3=2.337e-026 dpua1_4=5.6055e-042 dpua1_5=8.1436e-029 dketa_1=-0.0028179 dketa_2=0.00087739 dketa_3=0.0014002 dketa_4=2.8738e-018 dketa_5=0.00026796 dpketa_1=-1.0784e-017 dpketa_2=3.9912e-018 dpketa_3=-1.8696e-017 dpketa_4=-9.5866e-033 dpketa_5=-6.5149e-020 ss_flag_1=0.053919 ss_flag_2=-0.019956 ss_flag_3=0.093479 ss_flag_4=-9.5952e-017 ss_flag_5=0.00032575 ff_flag_1=-0.040011 ff_flag_2=0.0092905 ff_flag_3=0.14015 ff_flag_4=-7.6137e-017 ff_flag_5=0.0092578 monte_flag_1=0.0756092 monte_flag_2=-0.189108 monte_flag_3=-0.0582925 monte_flag_4=-0.707108 monte_flag_5=0.014055 sigma_local=1                          a_1=0.901479 b_1=0.000289007                c_1=0.00481065                 d_1=4.96369e-005 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1.07088                    b_2=-0.00531461                c_2=-0.010276 d_2=-0.000296336               a_3=0.972501                   b_3=-0.00703771 c_3=-0.00751154                d_3=-10.40812e-005             e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.69 b_4=0.0018                     c_4=0.011                      d_4=-0.00032 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=0.69                       b_5=-0.0012                    c_5=-0.006 d_5=0.00038                    e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=-0.0018                    mis_a_2=-0.086                     mis_a_3=0.14 mis_b_1=0.0019                     mis_b_2=-0.1555                    mis_b_3=0.1417 mis_c_1=0.1000                     mis_c_2=0.0000                     mis_c_3=0.0000 mis_d_1=0.00076                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.0024                     mis_e_2=-0.084                     mis_e_3=-0.063 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-3e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=60                         co_rsd=16.7 cf0=9e-011                     cco=0.92e-10 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.85                       l_rjtsswg=0                          ll_rjtsswg=0.0 w_rjtsswg=0.95                       ww_rjtsswg=1.0                        p_rjtsswg=0.0 noimod=6                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718                      tnoiamax=12117167.5188 tnoiac1=797021.1169                tnoiac2=8427254.9408               rnoiamax=0.4159 rnoiac1=0.013311                   rnoiac2=0.35427 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6               sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=1                   lreflod=0.9e-6              llodref=2 lod_clamp=-1e90 wlod0=0 ku00=-0e-9       lku00=0e-7        wku00=0e-8         pku00=0e-14 tku00=0           llodku00=1           wlodku00=1            kvsat0=0.5 kvth00=-3.8e-9     lkvth00=1.75e-8     wkvth00=3e-8         pkvth00=0e-15 llodvth0=1           wlodvth0=1 stk20=0           lodk20=1           steta00=5e-11        lodeta00=1 wlod00=0 ku000=0           lku000=-13e-32     wku000=0            pku000=0 llodku000=3           wlodku000=1 kvth000=0           lkvth000=3e-17       wkvth000=0            pkvth000=0e-14 llodvth00=1           wlodvth00=1 steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0           llod1=0.00e-6 ku01=2e-8        lku01=-3e-2       wku01=-5e-15     pku01=0 llodku01=-1          wlodku01=1           kvsat1=-0 kvth01=11e-9     lkvth01=-3e-24      wkvth01='1.5e-19'     pkvth01=0e-24 llodvth1=2           wlodvth1=1.5 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.1        lku02=0.4e-7      wku02=0            pku02=0 tku02=0           llodku02=1           wlodku02=1            kvsat2='0.4*0+0.5' kvth02=-0e-3       lkvth02=0e-8        wkvth02=0e-8         pkvth02=0 llodvth2=1           wlodvth2=1 stk22=0           lodk22=1           steta02=-1e-4        lodeta02=1 wlod02=0 ku002=0           lku002='-1.2e11*2'     wku002=3.5e-9       pku002=0 llodku002=-2          wlodku002=1 kvth002=0           lkvth002=-0e-11      wkvth002=0            pkvth002=0 llodvth02=1           wlodvth02=1 steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0.085        lku03=-0.05e-7        wku03=0e-7         pku03=0 tku03=0           llodku03=1           wlodku03=1            kvsat3=0.4 kvth03=0.1e-3      lkvth03=0e-20       wkvth03=0e-8         pkvth03=0e-20 llodvth3=3           wlodvth3=1 stk23=0           lodk23=1           steta03=0e-3         lodeta03=1 wlod03=0 ku003=0           lku003='-1.25e5*8e-1'     wku003=1.5e-9            pku003=0 llodku003=-1          wlodku003=1 kvth003=0e-3        lkvth003=-5e-26      wkvth003=-2e-10       pkvth003=0e-32 llodvth03=3           wlodvth03=1 steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.7                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=-1.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=-0.000              wkvth0dpl=0                   wdplkvth0=1 lkvth0dpl=0.0e-9              ldplkvth0=1.0                 pkvth0dpl=0 ku0dpl=1               wku0dpl=0                   wdplku0=1 lku0dpl=-4e-8              ldplku0=1                 pku0dpl=0 keta0dpl=0.00                wketa0dpl=0                   wdplketa0=1 kvsatdpl=0                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=1 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=1.0e-6              wkvth0dpx=0                   wdpxkvth0=1 lkvth0dpx=0                   ldpxkvth0=1                   pkvth0dpx=0 ku0dpx=0                   wku0dpx=0                   wdpxku0=1 lku0dpx=0                   ldpxku0=1                   pku0dpx=0 keta0dpx=0                   wketa0dpx=0                   wdpxketa0=1 kvsatdpx=0                   wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0.02               wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-2             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='0.5'               wku0dps=0                   wdpsku0=1 lku0dps='2e-8-0.5e-8'        ldpsku0=1.0                 pku0dps=0 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0.7                 wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=1 ku0dps_b1=0                 ku0dps_b2=0.11 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=0.002               wkvth0dpa=-1.0e-9            wdpakvth0=1 lkvth0dpa=0.010e-7            ldpakvth0=1.0                pkvth0dpa=-3.0e-17 ku0dpa=-0.1               wku0dpa=-10e-9               wdpaku0=1 lku0dpa=-0e-9               ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=1 ku0dpa_b1=-0.1             ku0dpa_b2=0.00 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2=-0.01               wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0.5e-9              ldp2kvth0=1                   pkvth0dp2=0 ku0dp2=0.1                wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=-0.0e-8              ldp2ku0=1.0                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0.00                wdp2=0 kvth0dp2l=-0.018              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.6               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0e-8               ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0.2                wdp2l=0 kvth0dp2l_b1=0.00            kvth0dp2l_b2=-0.016           dp2lbinflg=1 ku0dp2l_b1=-0.00            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=-0.007              wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=-0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.2              wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=-10.0e-5            ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=0.017           kvth0dp2a_b2=-0.02           dp2abinflg=1 ku0dp2a_b1=-0.12                ku0dp2a_b2=0.08 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx=-0.023              wkvth0enx=-0.0e-9             wenxkvth0=1.0 lkvth0enx=-11.0e-9              lenxkvth0=1.0                 pkvth0enx=-0.85e-16 ku0enx=-2.0                wku0enx=-1.0e-8             wenxku0=1.0 lku0enx=0.4e-7              lenxku0=1.0                 pku0enx=-7.0e-16 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=1.0                 wka0enx=0                   wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx=0.5                 wenx=0                   ku0enx0=-0.20 eny0=0.08e-6 enyref=0.08e-6             enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0.010               wkvth0eny=5.0e-10             wenykvth0=1 lkvth0eny=1.0e-8              lenykvth0=1.0                 pkvth0eny=0 ku0eny=14.0                wku0eny=1.0e-8              wenyku0=1 ku0eny0=0.04                wku0eny0=-1.0e-7             weny0ku0=1 lku0eny=8.0e-6              lenyku0=1.0                 pku0eny=2.0e-16 keta0eny=0e-4                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny=0.8                 weny=0 kvth0eny1=-6e-4              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=3.0e-18 ku0eny1=-1.5e-3            wku0eny1=-1.0e-10           weny1ku0=1 lku0eny1=-0.6e-8            leny1ku0=1.0                pku0eny1=-5.5e-17 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1=1.0e-8             weny1ka0=1 lka0eny1=4.0e-9             leny1ka0=1.0                pka0eny1=3.0e-15 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=0.045               wkvth0rx=0.0e-6              wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0e-15 ku0rx=0.05                wku0rx=0.0e-4              wrxku0=1.0 lku0rx=0.0e-7              lrxku0=1.0                 pku0rx=0.0e-14 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.4                 wrx=0                   ku0rx0=0.35 ry_mode=0 ryref=1.8027e-5           ringymax=1.8047e-5           ringymin=0.117e-6 kvth0ry=-0.0025             wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry='1.0e-8*0'           lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry=-0.8                 wku0ry=-0.5e-8             wryku0=1.0 lku0ry=4.0e-7               lryku0=1.0                 pku0ry=-2.0e-16 keta0ry=0.00                 wketa0ry=0                   wryketa0=1 kvsatry=0.7                 wry=0 kvth0ry0='-0.01*0'            ku0ry0='-0.14*0' sfxref=9.0e-8            sfxmax=1.53e-6          minwodx=0 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=0.0 kvth0odx1a=-0.009            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.07              lku0odx1a=1.6e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.6 kvth0odx1b=0.0000            lkvth0odx1b=2.7e-11           lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=0.0011            lku0odx1b=1.1e-6            lodx1bku0=0.5 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6 sfymax=1.53e-6           minwody=0.0e-6            wody=5e-7 kvth0odya=40                lkvth0odya=1.0e-4            lodyakvth0=1.0 wkvth0odya=1.8e-7            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=1                 lku0odya=1.0e-6            lodyaku0=1.0 wku0odya=-0.0e-8           wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=-1.5e-2           wketa0ody=0                 wodyketa0=1 kvsatody=0.0 lrefody=1.0e-7            lodyref=1 kvth0odyb=-0.00             lkvth0odyb=7.0e-17           lodybkvth0=2.0 wkvth0odyb=9.0e-9            wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.50             lku0odyb=0.6e-10           lodybku0=1.2 wku0odyb=-0.9e-7           wodybku0=1.0               pku0odyb=-1.8e-16 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model pch_mac.1 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.36641013 lvth0=2.2112744e-010             wvth0=-2.0903369e-009            pvth0=-1.5232419e-015 k2=0.080588658                lk2=-5.1267544e-008            wk2=-3.1676963e-008 pk2=2.0974631e-014             cit=0.0009153705               lcit=-2.336159e-011 wcit=4.409493e-011              pcit=3.5182555e-017             voff=-0.10833086 lvoff=-3.9833558e-009            wvoff=-6.2191677e-009            pvoff=1.9401964e-015 eta0=0.01251                    weta0=-2.27406e-009              etab=-0.0016752407 wetab=-4.6829865e-009            u0=0.00905957                 wu0=1.8033296e-009 ua=4.6248293e-010             lua=-2.9534622e-016            wua=2.2070636e-016 pua=2.2156991e-023             ub=5.737952e-019              lub=3.2448271e-026 wub=1.3303581e-025             pub=-2.16828e-033              uc=5.2857847e-010 luc=-5.090365e-016             wuc=-3.8207057e-018            puc=3.437489e-023 vsat=119473.86                  wvsat=-0.019433207               a0=1.6817965 la0=-9.9058032e-008            wa0=2.3309103e-007             pa0=-3.6037473e-013 ags=1.3791706                  lags=-1.4033597e-008            wags=-4.5170826e-008 pags=3.9856626e-013             keta=-0.30247196                lketa=1.9498265e-007 wketa=1.9955298e-007             pketa=-1.586007e-013             pclm=0.24285 wpclm=-7.95921e-008              pdiblc2=0.00022281481              lpdiblc2=1.5941351e-009 aigbacc=0.01112525                 waigbacc=5.116635e-010              aigc=0.0060012012 laigc=4.9887719e-012             waigc=-1.8183245e-011            paigc=-7.7296997e-018 aigsd=0.0047591237               laigsd=6.6715328e-012             waigsd=1.8015051e-010 paigsd=-6.0444087e-018            bigsd=0.000107568                wbigsd=9.8239392e-011 tvoff=0.00361771                 ltvoff=-5.6157e-010               wtvoff=-7.91667e-010 ptvoff=3.17148e-016               kt1=-0.14516631                lkt1=2.8301876e-012 wkt1=1.3652066e-009             pkt1=-6.9331164e-018            kt2=-0.07422012 wkt2=-1.1097413e-009            ute=-0.7132354                 wute=-1.0565283e-007 ua1=7.4150694e-010             lua1=2.7670499e-017             wua1=4.9331634e-016 pua1=-1.040477e-022             ub1=4.5355337e-019             lub1=-3.5939388e-026 wub1=-1.0454962e-024            pub1=3.2560905e-032             uc1=8.4523538e-010 luc1=-4.0698269e-016            wuc1=-1.2087892e-017            puc1=1.0875477e-022 at=90000                      jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=0 pu0=0                          lvsat=0                          pvsat=0 lpclm=0                          ppclm=0                          lat=0 leta0=0                          peta0=0                          wat=0 pat=0                          u0_mcl=-3.85649e-05               wu0_mcl=5.80825e-11 ags_ss=-0.388711                  ags_ff=0.388711                   ags_sf=0.310969 ags_fs=-0.310969                  lags_ss=3.48674e-07                lags_ff=-3.48674e-07 lags_sf=-2.7894e-07                lags_fs=2.7894e-07                 wags_ss=4.2e-13 wags_ff=-4.2e-13                   wags_sf=-3.3e-13                   wags_fs=3.3e-13 pags_ss=-4.7e-19                   pags_ff=4.7e-19                    pags_sf=-2.3e-19 pags_fs=2.3e-19                    lu0_mcl=3.45927e-11                pu0_mcl=-5.21e-17 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.2 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.34924706 lvth0=-1.5174147e-008            wvth0=-1.5192731e-008            pvth0=1.0229605e-014 k2=0.024853203                lk2=-1.2728403e-009            wk2=-9.5034947e-009 pk2=1.0850301e-015             cit=0.00079381841              lcit=8.5670635e-011 wcit=3.3476696e-010             pcit=-2.2555026e-016            voff=-0.10015073 lvoff=-1.1320931e-008            wvoff=-8.7511803e-009            pvoff=4.2114117e-015 eta0=0.01251                    weta0=-2.27406e-009              etab=-0.0016752407 wetab=-4.6829865e-009            u0=0.0061258891               wu0=3.8069735e-009 ua=3.9799559e-010             lua=-2.3750107e-016            wua=4.195386e-016 pua=-1.5619552e-022            ub=-3.1397633e-019            lub=8.2877933e-025 wub=7.2605976e-025             pub=-5.3411077e-031            uc=-1.4940575e-010 luc=9.9115344e-017             wuc=9.4830534e-017             puc=-5.4115273e-023 vsat=119484.18                  wvsat=-0.019442559               a0=1.7015983 la0=-1.1682019e-007            wa0=-3.3692499e-007            pa0=1.5092963e-013 ags=0.2566984                  lags=9.9282398e-007             wags=6.7536739e-007 pags=-2.4775652e-013            keta=0.002065                   lketa=-7.8187005e-008 wketa=-3.373189e-008             pketa=5.0655823e-014             pclm=-0.56037622 wpclm=2.0661048e-007             pdiblc2=0.0022759877               lpdiblc2=-2.47561e-010 aigbacc=0.011011265                waigbacc=1.0199159e-009             aigc=0.0060365241 laigc=-2.6695838e-011            waigc=-5.8214183e-011            paigc=2.8178052e-017 aigsd=0.0047492849               laigsd=1.5496933e-011             waigsd=3.0599515e-010 paigsd=-1.1892705e-016            bigsd=0.00011995288              wbigsd=2.1841285e-010 tvoff=0.00368386                 ltvoff=-6.20904e-010              wtvoff=-9.9288e-010 ptvoff=4.97636e-016               kt1=-0.13685972                lkt1=-7.4481821e-009 wkt1=1.2414151e-009             pkt1=1.0410785e-016             kt2=-0.073638265 wkt2=-4.4438771e-009            ute=-0.44341726                wute=-2.5225541e-007 ua1=5.6477922e-010             lua1=1.8619526e-016             wua1=3.9178507e-016 pua1=-1.2974152e-023            ub1=1.5569554e-018             lub1=-1.025691e-024 wub1=-1.6059667e-024            pub1=5.353029e-031              uc1=4.076418e-010 luc1=-1.4461255e-017            wuc1=2.1758206e-016             puc1=-9.7259181e-023 at=89999.997                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=2.6315117e-009 pu0=-1.7972686e-015            lvsat=-9.2589452e-006            pvsat=8.3886044e-012 lpclm=7.2049392e-007             ppclm=-2.5672371e-013            wpdiblc2=-4.1563753e-010 ppdiblc2=3.7282686e-016             laigbacc=1.0224454e-010             paigbacc=-4.5590241e-016 lbigsd=-1.1109237e-011            pbigsd=-1.0779559e-016            lkt2=-5.2192387e-010 pkt2=2.9907198e-015             lute=-2.4202687e-007            pute=1.3150252e-013 lat=2.6730599e-009             leta0=0                          peta0=0 wat=0                          pat=0                          ags_ss=-0.0794663 ags_ff=0.198666                   ags_sf=0.0993337                  ags_fs=-0.0993337 lags_ss=7.12817e-08                lags_ff=-1.78204e-07               lags_sf=-8.91024e-08 lags_fs=8.91024e-08                wags_ss=1.5e-13                    wags_ff=-3.7e-13 wags_sf=3.1e-13                    wags_fs=-3.1e-13                   pags_ss=3.9e-19 pags_ff=4e-20                      pags_sf=2e-20                      pags_fs=-2e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.3 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.37966145 lvth0=-1.5789153e-009            wvth0=5.6070339e-009             pvth0=9.3211045e-016 k2=0.028731632                lk2=-3.006498e-009             wk2=-6.6494526e-009 pk2=-1.9072673e-016            cit=0.00026012909              lcit=3.2422976e-010 wcit=-1.2783029e-009            pcit=4.9549198e-016             voff=-0.11927638 lvoff=-2.7717661e-009            wvoff=-2.6001223e-009            pvoff=1.4618888e-015 eta0=0.01251                    weta0=-2.27406e-009              etab=-0.0016752407 wetab=-4.6829865e-009            u0=0.010704245                wu0=4.1124742e-010 ua=7.2038608e-010             lua=-3.8160962e-016            wua=1.3025902e-016 pua=-2.6887552e-023            ub=1.3796263e-018             lub=7.1738953e-026 wub=-6.5430678e-025            pub=8.2913076e-032             uc=9.0618123e-011 luc=-8.1753264e-018            wuc=-4.3026067e-017            puc=7.5066279e-024 vsat=93905.876                  wvsat=0.016495591                a0=2.0740183 la0=-2.8329196e-007            wa0=9.537207e-007              pa0=-4.2598899e-013 ags=2.9126845                  lags=-1.9440179e-007            wags=2.3133634e-007 pags=-4.9274641e-014            keta=-0.12864799                lketa=-1.9758297e-008 wketa=4.5965312e-008             pketa=1.5031174e-014             pclm=1.1814019 wpclm=-5.4095381e-007            pdiblc2=0.0002230041               lpdiblc2=6.7012269e-010 aigbacc=0.01124                    aigc=0.0059352281               laigc=1.8583474e-011 waigc=3.1153831e-011             paigc=-1.1769451e-017            aigsd=0.0047366655 laigsd=2.11378e-011               waigsd=-4.7943902e-012            paigsd=1.9995875e-017 bigsd=2.4373077e-005             wbigsd=-4.3440377e-011            tvoff=0.00317943 ltvoff=-3.95423e-010              wtvoff=3.56139e-010               ptvoff=-1.05376e-016 kt1=-0.1333745                 lkt1=-9.0060768e-009            wkt1=2.0561997e-008 pkt1=-8.5321922e-015            kt2=-0.076087384               wkt2=2.733216e-009 ute=-0.96652301                wute=1.4051067e-008             ua1=2.3552202e-009 lua1=-6.1413184e-016            wua1=-8.0514659e-016            pua1=5.220543e-022 ub1=-3.5847646e-018            lub1=1.2726578e-024             wub1=1.5929991e-024 pub1=-8.9463481e-031            uc1=3.1544546e-010             luc1=2.6750507e-017 wuc1=1.2620654e-016             puc1=-5.6414323e-023            at=126410.26 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=5.8498672e-010             pu0=-2.7937905e-016            lvsat=0.011424242 pvsat=-1.6055964e-008            lpclm=-5.8080881e-008            ppclm=7.7437522e-014 wpdiblc2=2.6871226e-009             ppdiblc2=-1.0141069e-015            lbigsd=3.1614935e-011 pbigsd=9.2528003e-018             lkt2=5.7283251e-010             pkt2=-2.1744081e-016 lute=-8.1986029e-009            pute=1.2463522e-014             lat=-0.016275385 leta0=0                          peta0=0                          wat=0 pat=0                          vsat_ss=-7282.03                   vsat_ff=15527.6 vsat_sf=5461.55                    vsat_fs=-5461.55                   wvsat_ss=3.9e-08 wvsat_ff=-0.0124187                 wvsat_sf=2.1e-08                    wvsat_fs=-2.1e-08 ags_ss=-0.302311                  ags_ff=0.210505                   ags_sf=0.173078 ags_fs=-0.173078                  lags_ss=1.70891e-07                lags_ff=-1.83495e-07 lags_sf=-1.22066e-07               lags_fs=1.22066e-07                wags_ss=5.18e-12 wags_ff=-2.06982e-07               wags_sf=-2.2e-13                   wags_fs=2.2e-13 pags_ss=-3.82e-19                  pags_ff=9.25191e-14                pags_sf=1.27e-19 pags_fs=-1.27e-19                  lvsat_ss=0.00325507                 lvsat_ff=-0.00694083 lvsat_sf=-0.00244131                lvsat_fs=0.00244131                 pvsat_ss=-1.8e-15 pvsat_ff=5.55113e-09                pvsat_sf=-3.6e-15                   pvsat_fs=3.6e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.4 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.38281566 lvth0=-9.0706755e-010            wvth0=8.9973478e-009             pvth0=2.099736e-016 k2=0.026892186                lk2=-2.6146959e-009            wk2=-4.5495921e-009 pk2=-6.3799701e-016            cit=0.0015784893               lcit=4.3419033e-011 wcit=1.7069628e-009             pcit=-1.4036962e-016            voff=-0.11771705 lvoff=-3.1039026e-009            wvoff=7.3892067e-009             pvoff=-6.658383e-016 eta0=0.011213645                weta0=-1.0995621e-009            etab=-0.0016752523 wetab=-4.6829691e-009            u0=0.01146781                 wu0=2.3494676e-010 ua=-9.5928858e-010            lua=-2.3838913e-017            wua=1.3000123e-016 pua=-2.6832643e-023            ub=1.8440206e-018             lub=-2.717703e-026 wub=-3.8446608e-025            pub=2.5437006e-032             uc=4.5999857e-011 luc=1.3283642e-018             wuc=1.135589e-017              puc=-4.076729e-024 vsat=184431.28                  wvsat=-0.097940094               a0=2.7820758 la0=-4.3410821e-007            wa0=-1.7020677e-006            pa0=1.3969394e-013 ags=2.3646543                  lags=-7.7671363e-008            wags=2.9519465e-007 pags=-6.287646e-014             keta=-0.070121513               lketa=-3.2224437e-008 wketa=9.2308222e-008             pketa=5.1601342e-015             pclm=1.1347424 wpclm=-4.6340097e-007            pdiblc2=0.0043144648               lpdiblc2=-2.0135843e-010 aigbacc=0.010953218                waigbacc=6.8145998e-010             aigc=0.0060152241 laigc=1.5443185e-012             waigc=5.4077526e-013             paigc=-5.24887e-018 aigsd=0.0047298563               laigsd=2.2588167e-011             waigsd=9.9835281e-011 paigsd=-2.2902449e-018            bigsd=0.0001728                  tvoff=0.000778071 ltvoff=1.16066e-010               wtvoff=1.20844e-010               ptvoff=-5.52579e-017 kt1=-0.19799898                lkt1=4.7589377e-009             wkt1=-7.8829346e-009 pkt1=-2.4734218e-015            kt2=-0.078753557               wkt2=6.1528483e-009 ute=-0.84377831                wute=5.5465948e-008             ua1=-5.7361649e-010 lua1=9.7103693e-018             wua1=2.4471573e-015             pua1=-1.7068642e-022 ub1=3.2399604e-018             lub1=-1.8100859e-025            wub1=-4.0303232e-024 pub1=3.0313284e-031             uc1=4.6362342e-010             luc1=-4.8113977e-018 wuc1=-1.8413768e-016            puc1=9.6889949e-024             at=65003.033 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=4.2234741e-010             pu0=-2.4182701e-016            lvsat=-0.0078576689 pvsat=8.3188365e-009             lpclm=-4.8142427e-008            ppclm=6.0918768e-014 wpdiblc2=-3.5059508e-009            ppdiblc2=3.0501772e-016             laigbacc=6.1084647e-011 paigbacc=-1.4515098e-016            lkt2=1.1407272e-009             pkt2=-9.4582249e-016 lute=-3.4343223e-008            pute=3.6421524e-015             lat=-0.0031956455 leta0=2.7612367e-010             peta0=-2.5016804e-016            letab=2.4650642e-015 petab=-3.7123867e-021            wat=-0.014903579               pat=3.1744624e-009 vsat_ss=16285.8                    vsat_ff=-32289.3                   vsat_sf=-10142.8 vsat_fs=11523.8                    wvsat_ss=-2.9e-08                   wvsat_ff=0.0230632 wvsat_sf=4.7e-08                    wvsat_fs=5.3e-08                    ags_ss=0.845233 ags_ff=-1.10045                   ags_sf=-0.676192                  ags_fs=0.676192 lags_ss=-7.35356e-08               lags_ff=9.57397e-08                lags_sf=5.88287e-08 lags_fs=-5.88287e-08               wags_ss=-5e-13                     wags_ff=3.84386e-07 wags_sf=-3.6e-12                   wags_fs=3.6e-12                    pags_ss=1.4e-19 pags_ff=-3.34417e-14               pags_sf=2.9e-19                    pags_fs=-2.9e-19 pdiblc2_ss=0.00103571                 pdiblc2_fs=-0.00103571                lpdiblc2_ss=-2.20607e-10 lpdiblc2_fs=2.20607e-10                lvsat_ss=-0.00176486                lvsat_ff=0.00324417 lvsat_sf=0.000882425                lvsat_fs=-0.00117657                pvsat_ss=-5.8e-15 pvsat_ff=-2.0065e-09                pvsat_sf=4.3e-15                    pvsat_fs=-4.3e-15 wpdiblc2_ss=3e-16                      wpdiblc2_fs=-3e-16                     ppdiblc2_ss=4.1e-22 ppdiblc2_fs=-4.1e-22 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.5 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.42282363 lvth0=2.5736259e-009             wvth0=2.4136781e-008             pvth0=-1.1071571e-015 k2=0.070153724                lk2=-6.3784498e-009            wk2=-3.8797725e-008 pk2=2.3415906e-015             cit=-0.00045341499             lcit=2.2019471e-010 wcit=4.6202473e-010             pcit=-3.2060007e-017            voff=-0.14128279 lvoff=-1.0536837e-009            wvoff=6.9487028e-009             pvoff=-6.2751446e-016 eta0=0.014962618                weta0=-7.5123572e-009            etab=0.0079733369 wetab=-1.2245648e-008            u0=0.021631681                wu0=-7.218401e-009 ua=-8.3329164e-010            lua=-3.4800647e-017            wua=-6.5538895e-016 pua=4.1496303e-023             ub=1.6243584e-018             lub=-8.0664166e-027 wub=1.2341305e-026             pub=-9.085236e-033             uc=1.5384533e-010 luc=-8.0541917e-018            wuc=-1.1157175e-016            puc=6.6179757e-024 vsat=94326.615                  wvsat=-0.027184831               a0=-4.0096738 la0=1.5677401e-007             wa0=3.9217141e-006             pa0=-3.4957507e-013 ags=2.1403767                  lags=-5.815921e-008             wags=-1.0331813e-006 pags=5.2692244e-014             keta=-0.96541918                lketa=4.566646e-008 wketa=5.3284235e-007             pketa=-3.3166335e-014            pclm=0.33439753 wpclm=6.43455e-007               pdiblc2=0.00058333333              ppdiblc2=0 wpdiblc2=0                          lpdiblc2=1.2325e-010                aigbacc=0.011522839 waigbacc=-1.2994358e-009            aigc=0.006161488                laigc=-1.1180637e-011 waigc=-1.1037855e-010            paigc=4.4011113e-018             aigsd=0.0048384269 laigsd=1.3142521e-011             waigsd=1.5570334e-010             paigsd=-7.1507664e-018 bigsd=0.0001728                  tvoff=0.00287377                 ltvoff=-6.626e-011 wtvoff=-1.61564e-009              ptvoff=9.58163e-017               kt1=-0.093407899 lkt1=-4.3404865e-009            wkt1=-9.5906723e-008            pkt1=5.1846478e-015 kt2=-0.069475632               wkt2=-1.7679111e-008            ute=-1.2911104 wute=2.4777779e-007             ua1=6.3602592e-010             lua1=-9.5528521e-017 wua1=-4.5684023e-016            pua1=8.1961361e-023             ub1=-1.4038288e-018 lub1=2.2300107e-025             wub1=2.0675512e-024             pub1=-2.2738223e-031 uc1=3.4542e-010                luc1=5.4723e-018                wuc1=5.609348e-017 puc1=-1.1211116e-023            at=18565.371                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-4.6190937e-010 pu0=4.0661425e-016             lvsat=-1.8563051e-005            pvsat=2.1631286e-009 lpclm=2.1487581e-008             ppclm=-3.5377702e-014            laigbacc=1.1527573e-011 paigbacc=2.7186956e-017             lkt2=3.3354778e-010             pkt2=1.127558e-015 lute=4.5746703e-009             pute=-1.3088978e-014            lat=0.00084443108 leta0=-5.0037035e-011            peta0=3.0774513e-016             letab=-8.3942479e-010 petab=6.5794933e-016             wat=0.029020793                pat=-6.4695798e-010 vsat_ss=-8249.97                   vsat_ff=9250.01                    vsat_fs=-4833.28 wvsat_ss=2.4e-08                    wvsat_ff=-3e-08                     wvsat_fs=1.2e-08 a0_ss=-0.850004                  a0_fs=0.850004                   la0_ss=7.39501e-08 la0_fs=-7.39501e-08               wa0_ss=2.8e-12                    wa0_fs=-2.8e-12 pa0_ss=-1.2e-19                   pa0_fs=1.2e-19                    pdiblc2_ss=-0.0015 pdiblc2_fs=0.0015                     ppdiblc2_ss=7e-22                      ppdiblc2_fs=-7e-22 wpdiblc2_ss=-1.1e-15                   wpdiblc2_fs=1.1e-15                    lpdiblc2_ss=2.7e-16 lpdiblc2_fs=-2.7e-16                   ua1_ss=1.06664e-10                ua1_fs=1.77774e-10 lua1_ss=-9.27979e-18               lua1_fs=-1.54663e-17               wua1_ss=-9.66379e-17 wua1_fs=-1.61063e-16               pua1_ss=8.40749e-24                pua1_fs=1.40125e-23 lvsat_ss=0.000369754                lvsat_ff=-0.000369748               lvsat_fs=0.0002465 pvsat_ss=-8e-16                     pvsat_ff=1e-15                      pvsat_fs=-4.1e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.6 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.43718932 lvth0=3.3062759e-009             wvth0=8.5992859e-008             pvth0=-4.2618171e-015 k2=0.098710542                lk2=-7.8348475e-009            wk2=-2.6797381e-009 pk2=4.9957323e-016             cit=-0.0016801875              lcit=2.827601e-010 wcit=1.3016874e-009             pcit=-7.4882802e-017            voff=-0.18093686 lvoff=9.6867418e-010             wvoff=8.9393152e-008             pvoff=-4.8321813e-015 eta0=0.006317603                weta0=-2.0435871e-010            etab=-0.037622774 wetab=3.3382629e-009             u0=0.022530739                wu0=-8.7183962e-009 ua=-1.8100646e-009            lua=1.5014774e-017             wua=9.8659752e-017 pua=3.039819e-024              ub=2.4629583e-018             lub=-5.0835012e-026 wub=-6.6729713e-025            pub=2.5576324e-032             uc=1.0792e-010 luc=-5.712e-018                wuc=1.819248e-017              puc=-2.271587e-038 vsat=109693.84                  wvsat=-0.014207439               a0=14.661101 la0=-7.954355e-007             wa0=-3.3657071e-006            pa0=2.2083407e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.48706011                lketa=2.1270147e-008 wketa=-3.7602142e-008            pketa=-4.0736657e-015            pclm=0.58307469 wpclm=9.600641e-008              pdiblc2=0.003                      ppdiblc2=0 wpdiblc2=0                          lpdiblc2=0                          aigbacc=0.014123597 waigbacc=-4.3426966e-009            aigc=0.0062078342               laigc=-1.3544298e-011 waigc=-1.3979845e-010            paigc=5.9015259e-018             aigsd=0.0050135744 laigsd=4.2099999e-012             waigsd=5.4439624e-011             paigsd=-1.9863167e-018 bigsd=0.0001728                  tvoff=0.00318342                 ltvoff=-8.2052e-011 wtvoff=-9.11379e-010              ptvoff=5.9899e-017                kt1=-0.14551862 lkt1=-1.68284e-009              wkt1=-3.5061027e-008            pkt1=2.0815173e-015 kt2=-0.14452781                wkt2=5.2790029e-008             ute=-0.34968367 wute=-1.3491998e-006            ua1=4.8034798e-010             lua1=-8.7588946e-017 wua1=-2.6190285e-016            pua1=7.2019555e-023             ub1=3.6729192e-018 lub1=-3.5913077e-026            wub1=-3.2537592e-024            pub1=4.40046e-032 uc1=1.5549807e-009             luc1=-5.6215298e-017            wuc1=-9.9326055e-016 puc1=4.230594e-023              at=-64019.03                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-5.0776135e-010 pu0=4.83114e-016               lvsat=-0.0008022917              pvsat=1.5012816e-009 lpclm=8.8050457e-009             ppclm=-7.4578237e-015            laigbacc=-1.2111106e-010 paigbacc=1.8239326e-016             lkt2=4.1612087e-009             pkt2=-2.4663682e-015 lute=-4.3438094e-008            pute=6.8356879e-014             lat=0.0050562355 leta0=3.9085875e-010             peta0=-6.4962795e-017            letab=1.4859769e-009 petab=-1.3683011e-016            wat=0.064787015                pat=-2.4710353e-009 u0_ss=0.00234243                 u0_ff=-0.00234243                wu0_ss=-2.12224e-09 wu0_ff=2.12224e-09                vsat_ss=-999.959                   vsat_ff=6666.62 wvsat_ss=5.2e-08                    wvsat_ff=-4e-09                     a0_ss=0.599996 a0_ff=-2.11365                   a0_sf=2.11365                    a0_fs=-0.599996 la0_ss=7e-14                      la0_ff=1.07796e-07                la0_sf=-1.07796e-07 la0_fs=-7e-14                     wa0_ss=-1.1e-12                   wa0_ff=3.18336e-06 wa0_sf=-3.18336e-06               wa0_fs=1.1e-12                    pa0_ss=-2.1e-19 pa0_ff=-1.62352e-13               pa0_sf=1.62352e-13                pa0_fs=2.1e-19 pdiblc2_ss=-0.00150004                pdiblc2_fs=0.00150004                 ppdiblc2_ss=3e-23 ppdiblc2_fs=-3e-23                     wpdiblc2_ss=2.8e-14                    wpdiblc2_fs=-2.8e-14 lpdiblc2_ss=-1.7e-16                   lpdiblc2_fs=1.7e-16                    ua1_ss=-7.52922e-11 ua1_fs=-1.25487e-10               lua1_ss=3e-24                      lua1_fs=6e-24 wua1_ss=6.82154e-17                wua1_fs=1.13691e-16                pua1_ss=3.9e-29 pua1_fs=-1e-30                     lu0_ss=-1.19464e-10               lu0_ff=1.19464e-10 pu0_ss=1.08234e-16                pu0_ff=-1.08234e-16               lvsat_ss=-1.1e-10 lvsat_ff=-0.000238                  pvsat_ss=2e-17                      pvsat_ff=-4e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.7 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.25564864 lvth0=-4.3184327e-009            wvth0=-2.0712982e-007            pvth0=8.0493354e-015 k2=0.046671069                lk2=-5.6491896e-009            wk2=1.3026108e-008 pk2=-1.600723e-016             cit=-0.0024617377              lcit=3.1558521e-010 wcit=-8.5527514e-009            pcit=3.3900363e-016             voff=0.0021579669 lvoff=-6.7213086e-009            wvoff=-1.5857707e-007            pvoff=5.5825682e-015 eta0=0.0073469933               weta0=-5.0189696e-009            etab=-0.018088644 wetab=3.4256689e-009             u0=0.0064544946               wu0=1.2395451e-008 ua=-8.192925e-010             lua=-2.6597654e-017            wua=-5.8341867e-016 pua=3.1687113e-023             ub=2.5043231e-019             lub=4.2091079e-026 wub=1.3962028e-024             pub=-6.1090671e-032            uc=-3.9886507e-012 luc=-1.0118367e-018            wuc=3.6229718e-017             puc=-7.5756397e-025 vsat=57938.424                  wvsat=0.0043888774               a0=30.786936 la0=-1.4727206e-006            wa0=-3.4462703e-005            pa0=1.3281572e-012 ags=1                          lags=0                          wags=0 pags=0                          keta=0.7162087                  lketa=-2.9267143e-008 wketa=-1.1950866e-006            pketa=4.4540681e-014             pclm=0.92602378 wpclm=2.4938649e-007             pdiblc2=-0.0025366667              lpdiblc2=2.3254e-010 aigbacc=0.0068826433               waigbacc=6.5621791e-009             aigc=0.0063251189 laigc=-1.8470253e-011            waigc=-4.4994445e-010            paigc=1.8927658e-017 aigsd=0.0024382071               laigsd=1.1237543e-010             waigsd=2.4312454e-009 paigsd=-1.0181216e-016            bigsd=-0.0026436041              wbigsd=2.5516621e-009 tvoff=-0.0010626                 ltvoff=9.62804e-011               wtvoff=4.32439e-009 ptvoff=-1.60003e-016              kt1=-0.29478664                lkt1=4.5864171e-009 wkt1=3.117102e-007              pkt1=-1.2482874e-014            kt2=-0.067960279 wkt2=-7.4651871e-009            ute=-1.3715087                 wute=2.0663625e-007 ua1=-2.0823689e-009            lua1=2.0045163e-017             wua1=1.8252017e-015 pua1=-1.5638835e-023            ub1=5.4443821e-018             lub1=-1.1031452e-025 wub1=-4.8383688e-024            pub1=1.105582e-031              uc1=3.4854687e-010 luc1=-5.5450752e-018            wuc1=5.3906062e-017             puc1=-1.6750579e-024 at=69499.318                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=1.6744092e-010 pu0=-4.0366757e-016            lvsat=0.0013714359               pvsat=7.202363e-010 lpclm=-5.5988158e-009            ppclm=-1.3899787e-014            wpdiblc2=8.33822e-009 ppdiblc2=-3.5020524e-016            laigbacc=1.8300898e-010             paigbacc=-2.7561152e-016 lbigsd=1.1828897e-010             pbigsd=-1.0716981e-016            lkt2=9.453725e-010 pkt2=6.4350913e-017             lute=-5.21444e-010              pute=3.0117651e-015 lat=-0.00055153513             leta0=3.4762435e-010             peta0=1.3725086e-016 letab=6.6554341e-010             petab=-1.4050116e-016            wat=-0.08087985 pat=3.646973e-009              cit_mc=0.00553574                 lcit_mc=-2.32501e-10 wcit_mc=-8.33738e-09               pcit_mc=3.5017e-16                 voff_ss=-0.0110715 voff_sf=0.00733331                 voff_mc=0.0664289                  lvoff_ss=4.65003e-10 lvoff_sf=-3.08001e-10               lvoff_mc=-2.79002e-09               wvoff_ss=1.66748e-08 wvoff_sf=-3.2e-14                   wvoff_mc=-1.00049e-07               pvoff_ss=-7.0034e-16 pvoff_sf=-2.6e-22                   pvoff_mc=4.20204e-15                eta0_mc=0.00664289 eta0_mcl=0.0127322                  weta0_mc=-1.00049e-08               weta0_mcl=-1.9176e-08 u0_ss=-0.00455673                u0_ff=0.00344958                 u0_sf=0.000830362 u0_fs=-0.00110715                wu0_ss=5.45719e-09                wu0_ff=-3.78972e-09 wu0_sf=-1.25061e-09               wu0_fs=1.66748e-09                vsat_ss=6404.83 vsat_ff=-6404.83                   vsat_mc=-33214.5                   vsat_mcl=-38750.2 wvsat_ss=-0.0166748                 wvsat_ff=0.0166748                  wvsat_mc=0.0500243 wvsat_mcl=0.0583617                  a0_ss=2.8                        a0_ff=2.11365 a0_sf=-2.11365                   a0_fs=-2.8                       la0_ss=-9.24002e-08 la0_ff=-6.97504e-08               la0_sf=6.97504e-08                la0_fs=9.24002e-08 wa0_ss=-3e-13                     wa0_ff=-3.18336e-06               wa0_sf=3.18336e-06 wa0_fs=3e-13                      pa0_ss=-8e-20                     pa0_ff=1.05051e-13 pa0_sf=-1.05051e-13               pa0_fs=8e-20                      pdiblc2_ss=-0.00699996 pdiblc2_fs=0.00699996                 lpdiblc2_ss=2.31e-10                   lpdiblc2_fs=-2.31e-10 ua1_ss=-6.27437e-10               ua1_fs=-1.04573e-09               lua1_ss=2.319e-17 lua1_fs=3.86502e-17                wua1_ss=5.68458e-16                wua1_fs=9.4743e-16 pua1_ss=-2.10102e-23               pua1_fs=-3.5017e-23                lu0_ss=1.70301e-10 lu0_ff=-1.23801e-10               lu0_sf=-3.48752e-11               lu0_fs=4.65003e-11 pu0_ss=-2.10102e-16               pu0_ff=1.40068e-16                pu0_sf=5.25255e-17 pu0_fs=-7.0034e-17                lvsat_ss=-0.000311003               lvsat_ff=0.000311003 lvsat_mc=0.00139501                 lvsat_mcl=0.00162751                 pvsat_ss=7.0034e-10 pvsat_ff=-7.0034e-10                pvsat_mc=-2.10102e-09               pvsat_mcl=-2.45119e-09 wpdiblc2_ss=-2.4e-14                   wpdiblc2_fs=2.4e-14                    ppdiblc2_ss=2e-22 ppdiblc2_fs=-2e-22                     leta0_mc=-2.79002e-10               leta0_mcl=-5.34753e-10 peta0_mc=4.20204e-16                peta0_mcl=8.05391e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_mac.8 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.36832197 lvth0=-6.4493279e-009            wvth0=-3.5821282e-010            pvth0=4.5201907e-015 k2=0.065956963                lk2=-4.1033462e-008            wk2=-1.8420646e-008 pk2=1.1702553e-014             cit=0.0013283504               lcit=3.8936065e-011 wcit=-3.3006486e-010            pcit=-2.1259121e-017            voff=-0.10871167 lvoff=-4.6379088e-009            wvoff=-5.8741499e-009            pvoff=2.5332214e-015 eta0=0.010025783                weta0=-2.33597e-011              etab=-0.0068119467 wetab=-2.913092e-011             u0=0.0111865                  wu0=-1.23669e-010 ua=1.2051206e-009             lua=-3.0863158e-016            wua=-4.5212338e-016 pua=3.4193533e-023             ub=1.7400376e-019             lub=4.5599575e-026 wub=4.9524685e-025             pub=-1.4083361e-032            uc=6.522513e-010 luc=-6.3924857e-016            wuc=-1.1586829e-016            puc=1.5234702e-022 vsat=86700.057                  wvsat=0.010259855                a0=2.1066518 la0=-7.2740885e-007            wa0=-1.5182789e-007            pa0=2.0891111e-013 ags=1.2786652                  lags=4.3195267e-007             wags=4.5887073e-008 pags=-5.4972951e-015            keta=-0.17786492                lketa=6.1763702e-008 wketa=8.6658997e-008             pketa=-3.7904334e-014            pclm=0.17775 wpclm=-2.0611502e-008            pdiblc2=0.00022281481              lpdiblc2=1.5941351e-009 aigbacc=0.011350267                waigbacc=3.077984e-010              aigc=0.0059775085 laigc=4.5449182e-012             waigc=3.2823156e-012             paigc=-7.3275683e-018 aigsd=0.0046286251               waigsd=2.9838226e-010             bigsd=-0.00011945633 wbigsd=3.0392344e-010             tvoff=0.00279636                 ltvoff=-4.89297e-010 wtvoff=-4.75267e-011              ptvoff=2.51668e-016               kt1=-0.15277318 lkt1=-1.7840448e-011            wkt1=8.2570301e-009             pkt1=1.1794479e-017 kt2=-0.0747079                 wkt2=-6.678126e-010             ute=-0.79766633 wute=-2.9158402e-008            ua1=1.7324235e-009             lua1=-2.199844e-016 wua1=-4.0445404e-016            pua1=1.2032764e-022             ub1=-1.1873031e-018 lub1=2.1497733e-026             wub1=4.411197e-025              pub1=-1.9477126e-032 uc1=8.4398622e-010             luc1=-3.9574404e-016            wuc1=-1.0956157e-017 puc1=9.8572547e-023             at=90000                      jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=0 pu0=0                          lvsat=0                          pvsat=0 lpclm=-1.5111072e-014            ppclm=1.3690632e-020             lat=0 leta0=0                          peta0=0                          wat=0 pat=0                          u0_mcl=6.42855e-05                wu0_mcl=-3.50999e-11 ags_ss=-0.388711                  ags_ff=0.388711                   ags_sf=0.310969 ags_fs=-0.310969                  lags_ss=3.48674e-07                lags_ff=-3.48674e-07 lags_sf=-2.78939e-07               lags_fs=2.78939e-07                wags_ss=-4.3e-13 wags_ff=4.3e-13                    wags_sf=-2.6e-13                   wags_fs=2.6e-13 pags_ss=2e-19                      pags_ff=-2e-19                     pags_sf=4.4e-19 pags_fs=-4.4e-19                   lu0_mcl=-5.76641e-11               pu0_mcl=3.14846e-17 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.9 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.36541853 lvth0=-9.0537129e-009            wvth0=-5.413798e-010             pvth0=4.6844914e-015 k2=0.019323197                lk2=7.9702636e-010             wk2=-4.4933087e-009 pk2=-7.9026908e-016            cit=0.0014269315               lcit=-4.9491184e-011 wcit=-2.388335e-010             pcit=-1.0309365e-016            voff=-0.10494878 lvoff=-8.0132265e-009            wvoff=-4.4041502e-009            pvoff=1.2146317e-015 eta0=0.010025783                weta0=-2.33597e-011              etab=-0.0068119467 wetab=-2.913092e-011             u0=0.011559613                wu0=-1.1159799e-009 ua=1.9267163e-009             lua=-9.5590294e-016            wua=-9.654824e-016 pua=4.9467658e-022             ub=-6.3969102e-019            lub=7.754838e-025 wub=1.0211573e-024             pub=-4.8582501e-031            uc=-1.9185533e-010 luc=1.1791508e-016             wuc=1.3328985e-016             puc=-7.1147832e-023 vsat=86700.057                  wvsat=0.010259855                a0=1.7736404 la0=-4.2869764e-007            wa0=-4.0219522e-007            pa0=4.334906e-013 ags=1.2063666                  lags=4.9680452e-007             wags=-1.85032e-007 pags=2.0163711e-013             keta=-0.10601775                lketa=-2.6832143e-009 wketa=6.4191078e-008             pketa=-1.7750611e-014            pclm=-0.31952263 wpclm=-1.1602873e-008            pdiblc2=0.0024793578               lpdiblc2=-4.2998398e-010 aigbacc=0.011459798                waigbacc=6.1354481e-010             aigc=0.0059933191 laigc=-9.6371856e-012            waigc=-1.9070506e-011            paigc=1.2722912e-017 aigsd=0.0045989734               laigsd=2.6597551e-011             waigsd=4.4217736e-010 paigsd=-1.2898421e-016            bigsd=-0.00015277571             wbigsd=4.6550496e-010 tvoff=0.00236575                 ltvoff=-1.03036e-010              wtvoff=2.01325e-010 ptvoff=2.84481e-017               kt1=-0.13444828                lkt1=-1.6455281e-008 wkt1=-9.4335408e-010            pkt1=8.2645391e-015             kt2=-0.073831813 wkt2=-4.2685226e-009            ute=-0.60845786                wute=-1.0272863e-007 ua1=1.1450799e-009             lua1=3.0686275e-016             wua1=-1.3396738e-016 pua1=-1.222989e-022             ub1=-4.484135e-019             lub1=-6.412862e-025 wub1=2.1089753e-025             pub1=1.8703216e-031             uc1=5.9993048e-010 luc1=-1.7682604e-016            wuc1=4.336852e-017              puc1=4.9843312e-023 at=89999.997                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-3.3468196e-010 pu0=8.9010287e-016             lvsat=0                          pvsat=0 lpclm=4.4605354e-007             ppclm=-8.0807261e-015            wpdiblc2=-5.9989084e-010 ppdiblc2=5.3810208e-016             laigbacc=-9.8249805e-011            paigbacc=-2.7425453e-016 lbigsd=2.9887484e-011             pbigsd=-1.4493862e-016            lkt2=-7.8584994e-010 pkt2=3.2298368e-015             lute=-1.6972001e-007            pute=6.5992496e-014 lat=2.67306e-009               leta0=0                          peta0=0 wat=0                          pat=0                          ags_ss=-0.0794666 ags_ff=0.198667                   ags_sf=0.0993334                  ags_fs=-0.0993334 lags_ss=7.12816e-08                lags_ff=-1.78204e-07               lags_sf=-8.9102e-08 lags_fs=8.9102e-08                 wags_ss=-1.5e-13                   wags_ff=-1.3e-13 wags_sf=-7e-14                     wags_fs=7e-14                      pags_ss=4.7e-20 pags_ff=-1.2e-19                   pags_sf=-6e-20                     pags_fs=6e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.10 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.38517628 lvth0=-2.2199781e-010            wvth0=1.0603471e-008             pvth0=-2.9725678e-016 k2=0.026414214                lk2=-2.3726584e-009            wk2=-4.5498718e-009 pk2=-7.6498537e-016            cit=0.00027395986              lcit=4.6588714e-010 wcit=-1.2908336e-009            pcit=3.6715039e-016             voff=-0.11719957 lvoff=-2.5371217e-009            wvoff=-4.48171e-009              pvoff=1.2493009e-015 eta0=0.010025783                weta0=-2.33597e-011              etab=-0.0068119467 wetab=-2.913092e-011             u0=0.010301312                wu0=7.763047e-010 ua=5.7184747e-010             lua=-3.5027656e-016            wua=2.64835e-016 pua=-5.52753e-023              ub=9.1332373e-019             lub=8.1286206e-026 wub=-2.3183664e-025            pub=7.4263265e-032             uc=9.8578554e-011 luc=-1.1908865e-017            wuc=-5.0238217e-017            puc=1.0889214e-023 vsat=107432.41                  wvsat=0.0042405538               a0=2.1520053 la0=-5.9782673e-007            wa0=8.830645e-007              pa0=-1.4102049e-013 ags=2.607053                   lags=-1.2930228e-007            wags=5.0823849e-007 pags=-1.082548e-013             keta=-0.05965975                lketa=-2.3405239e-008 wketa=-1.6538037e-008            pketa=1.8335304e-014             pclm=0.58987536 wpclm=-5.0308025e-009            pdiblc2=0.003185705                lpdiblc2=-7.4572117e-010 aigbacc=0.01124                    aigc=0.0059597305               laigc=5.3769095e-012 waigc=8.9545866e-012             paigc=1.9569623e-019             aigsd=0.0044675343 laigsd=8.5350828e-011             waigsd=2.3903848e-010             paigsd=-3.8181128e-017 bigsd=-0.0003214088              wbigsd=2.6983801e-010             tvoff=0.00321438 ltvoff=-4.82376e-010              wtvoff=3.24467e-010               ptvoff=-2.65965e-017 kt1=-0.15351877                lkt1=-7.9307689e-009            wkt1=3.8812709e-008 pkt1=-9.5064212e-015            kt2=-0.078819456               wkt2=5.2084732e-009 ute=-1.0387511                 wute=7.9489747e-008             ua1=2.2343177e-009 lua1=-1.8002653e-016            wua1=-6.9560896e-016            pua1=1.2875489e-022 ub1=-3.1229237e-018            lub1=5.5421987e-025             wub1=1.1745713e-024 pub1=-2.4373002e-031            uc1=2.1655592e-010             luc1=-5.4576112e-018 wuc1=2.1580047e-016             puc1=-2.7233768e-023            at=165635.3 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=2.2777843e-010             pu0=4.4251659e-017             lvsat=-0.0092673607 pvsat=2.6906277e-009             lpclm=3.9552633e-008             ppclm=-1.1018442e-014 wpdiblc2=2.9155583e-012             ppdiblc2=2.6864762e-016             lbigsd=1.0526648e-010 pbigsd=-5.7475495e-017            lkt2=1.4436266e-009             pkt2=-1.0063803e-015 lute=2.2621089e-008             pute=-1.5459119e-014            lat=-0.033808976 leta0=0                          peta0=0                          wat=-0.035537883 pat=1.5885434e-008             vsat_ss=-7282.06                   vsat_ff=1820.51 vsat_sf=5461.57                    vsat_fs=-5461.57                   wvsat_ss=3.3e-08 wvsat_ff=-3.3e-09                   wvsat_sf=0.0                        wvsat_fs=0.0 ags_ss=-0.302311                  ags_ff=-0.0179486                 ags_sf=0.173077 ags_fs=-0.173077                  lags_ss=1.70892e-07                lags_ff=-8.13771e-08 lags_sf=-1.22066e-07               lags_fs=1.22066e-07                wags_ss=6.7e-13 wags_ff=3.3e-13                    wags_sf=6.7e-13                    wags_fs=-6.7e-13 pags_ss=8.8e-20                    pags_ff=3e-20                      pags_sf=-8.5e-20 pags_fs=8.5e-20                    lvsat_ss=0.00325507                 lvsat_ff=-0.000813773 lvsat_sf=-0.00244131                lvsat_fs=0.00244131                 pvsat_ss=1.2e-15 pvsat_ff=-3e-16                     pvsat_sf=-9e-16                     pvsat_fs=9e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.11 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.38358961 lvth0=-5.599589e-010             wvth0=9.6985415e-009             pvth0=-1.0450684e-016 k2=0.030860038                lk2=-3.319619e-009             wk2=-8.1444665e-009 pk2=6.6328258e-019             cit=0.0025296214               lcit=-1.4568762e-011 wcit=8.4523716e-010             pcit=-8.7832677e-017            voff=-0.1139599 lvoff=-3.2271714e-009            wvoff=3.9852273e-009             pvoff=-5.5415675e-016 eta0=0.010025784                weta0=-2.335989e-011             etab=-0.0068119138 wetab=-2.9153786e-011            u0=0.011569345                wu0=1.4295543e-010 ua=-7.1976534e-010            lua=-7.5163032e-017            wua=-8.7006826e-017 pua=1.9667009e-023             ub=1.175205e-018              lub=2.5505504e-026 wub=2.2148089e-025             pub=-2.2293369e-032            uc=5.6699869e-011 luc=-2.9887056e-018            wuc=1.6616797e-018             puc=-1.6546374e-025 vsat=57019.093                  wvsat=0.017495347                a0=1.0978825 la0=-3.7329857e-007            wa0=-1.7618854e-007            pa0=8.4600408e-014 ags=2.6904762                  lags=-1.4707143e-007            wags=0 pags=0                          keta=-0.012400347               lketa=-3.3471492e-008 wketa=4.0012846e-008             pketa=6.2899655e-015             pclm=0.72561484 wpclm=-9.2731359e-008            pdiblc2=-0.0019140159              lpdiblc2=3.4051938e-010 aigbacc=0.011587045                waigbacc=1.0721252e-010             aigc=0.0060091669 laigc=-5.1530445e-012            waigc=6.0285556e-012             paigc=8.1894084e-019 aigsd=0.0047366147               laigsd=2.8036702e-011             waigsd=9.3712137e-011 paigsd=-7.2266172e-018            bigsd=0.0001728                  tvoff=0.000432603 ltvoff=1.10144e-010               wtvoff=4.33838e-010               ptvoff=-4.98926e-017 kt1=-0.18596507                lkt1=-1.0197087e-009            wkt1=-1.8785662e-008 pkt1=2.7620318e-015             kt2=-0.068514661               wkt2=-3.123591e-009 ute=-0.67795565                wute=-9.4769387e-008            ua1=2.6844185e-009 lua1=-2.7589801e-016            wua1=-5.0462248e-016            pua1=8.8074769e-023 ub1=-1.6965369e-018            lub1=2.5039947e-025             wub1=4.4214332e-025 pub1=-8.7722861e-032            uc1=1.0466984e-010             luc1=1.8374124e-017 wuc1=1.4107427e-016             puc1=-1.1317088e-023            at=-22583.277 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=-4.2312711e-011            pu0=1.7915505e-016             lvsat=0.0014706752 pvsat=-1.3264328e-010            lpclm=1.0640124e-008             ppclm=7.6617768e-015 wpdiblc2=2.1370527e-009             ppdiblc2=-1.8592358e-016            laigbacc=-7.3920551e-011 paigbacc=-2.2836266e-017            lkt2=-7.5129478e-010            pkt2=7.6834941e-016 lute=-5.4228349e-008            pute=2.1658076e-014             lat=0.0062815799 leta0=-4.4611667e-017            peta0=4.0418169e-023             letab=-7.0081987e-015 petab=4.8703895e-021             wat=0.064449617                pat=-5.4119038e-009 vsat_ss=16285.7                    vsat_ff=-6833.32                   vsat_sf=-10142.9 vsat_fs=11523.8                    wvsat_ss=-3.3e-08                   wvsat_ff=3.3e-09 wvsat_sf=0.0                        wvsat_fs=0.0                        ags_ss=0.845236 ags_ff=-0.676194                  ags_sf=-0.676194                  ags_fs=0.676194 lags_ss=-7.35358e-08               lags_ff=5.88287e-08                lags_sf=5.88287e-08 lags_fs=-5.88287e-08               wags_ss=1.7e-12                    wags_ff=-3.3e-13 wags_sf=-3.3e-13                   wags_fs=3.3e-13                    pags_ss=-4.3e-19 pags_ff=4e-20                      pags_sf=4e-20                      pags_fs=-4e-20 pdiblc2_ss=0.00103572                 pdiblc2_fs=-0.00103572                lpdiblc2_ss=-2.20607e-10 lpdiblc2_fs=2.20607e-10                lvsat_ss=-0.00176486                lvsat_ff=0.0010295 lvsat_sf=0.00088243                 lvsat_fs=-0.00117657                pvsat_ss=3.2e-15 pvsat_ff=4.7e-15                    pvsat_sf=-4.9e-15                   pvsat_fs=4.9e-15 wpdiblc2_ss=-5e-15                     wpdiblc2_fs=5e-15                      ppdiblc2_ss=-2.8e-22 ppdiblc2_fs=2.8e-22 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.12 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.42618247 lvth0=3.1456204e-009             wvth0=2.717989e-008              pvth0=-1.6253841e-015 k2=0.03967263                 lk2=-4.0863145e-009            wk2=-1.1181854e-008 pk2=2.6491601e-016             cit=-0.00036625196             lcit=2.3737222e-010 wcit=3.8305502e-010             pcit=-4.7622831e-017            voff=-0.13757322 lvoff=-1.1728129e-009            wvoff=3.5878321e-009             pvoff=-5.1958337e-016 eta0=0.0059811284               weta0=6.2487264e-010             etab=-0.0030104229 wetab=-2.2943615e-009            u0=0.011960667                wu0=1.543537e-009 ua=-1.8104847e-009            lua=1.9729557e-017             wua=2.2994801e-016 pua=-7.908062e-024             ub=1.8400964e-018             lub=-3.2340049e-026 wub=-1.8311732e-025            pub=1.2906675e-032             uc=4.8527306e-011 luc=-2.2776926e-018            wuc=-1.6153623e-017            puc=1.3844675e-024 vsat=30426.022                  wvsat=0.030709106                a0=-1.3915797 la0=-1.5671536e-007            wa0=1.5497208e-006             pa0=-6.5553703e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.605301                  lketa=1.8110865e-008 wketa=2.0657528e-007             pketa=-8.200966e-015             pclm=1.1595335 wpclm=-1.0411822e-007            pdiblc2=0.00058333333              ppdiblc2=0 wpdiblc2=0                          lpdiblc2=1.2325e-010                aigbacc=0.010019322 waigbacc=6.2750567e-011             aigc=0.0059956228               laigc=-3.9747039e-012 waigc=3.9895284e-011             paigc=-2.1274645e-018            aigsd=0.0050020492 laigsd=4.9438992e-012             waigsd=7.4615416e-012             paigsd=2.7718457e-019 bigsd=0.0001728                  tvoff=0.000876532                ltvoff=7.15219e-011 wtvoff=1.93855e-010               ptvoff=-2.90141e-017              kt1=-0.21957747 lkt1=1.9045705e-009             wkt1=1.840291e-008              pkt1=-4.7337392e-016 kt2=-0.094547962               wkt2=5.03642e-009               ute=-1.3158522 wute=2.7019386e-007             ua1=-1.5151623e-009            lua1=8.9465528e-017 wua1=1.4921363e-015             pua1=-8.5643247e-023            ub1=3.3153533e-018 lub1=-1.8563497e-025            wub1=-2.2080277e-024            pub1=1.4284202e-031 uc1=4.2957778e-010             luc1=-9.8928667e-018            wuc1=-2.0153467e-017 puc1=2.7097252e-024             at=43143.906                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-7.6357724e-011 pu0=5.7304456e-017             lvsat=0.0037842724               pvsat=-1.2822404e-009 lpclm=-2.7110803e-008            ppclm=8.652434e-015              laigbacc=6.2471317e-011 paigbacc=-1.8968076e-017            lkt2=1.5136024e-009             pkt2=5.842845e-017 lute=1.2686533e-009             pute=-1.0093726e-014            lat=0.00056331496 leta0=3.5188495e-010             peta0=-5.639619e-017             letab=-3.3073672e-010 petab=1.9707794e-016             wat=0.0067526396               pat=-3.9226678e-010 vsat_ss=-8249.99                   vsat_ff=9250.01                    vsat_fs=-4833.34 wvsat_ss=3.3e-08                    wvsat_ff=8e-09                      wvsat_fs=-3.3e-09 a0_ss=-0.850003                  a0_fs=0.850003                   la0_ss=7.39505e-08 la0_fs=-7.39505e-08               wa0_ss=5e-12                      wa0_fs=-5e-12 pa0_ss=-3e-19                     pa0_fs=3e-19                      pdiblc2_ss=-0.0015 pdiblc2_fs=0.0015                     ppdiblc2_ss=7.4e-22                    ppdiblc2_fs=-7.4e-22 wpdiblc2_ss=7.5e-15                    wpdiblc2_fs=-7.5e-15                   lpdiblc2_ss=2.5e-16 lpdiblc2_fs=-2.5e-16                   lvsat_ss=0.000369753                lvsat_ff=-0.000369754 lvsat_fs=0.0002465                  pvsat_ss=3e-16                      pvsat_ff=-1.3e-16 pvsat_fs=-3.5e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.13 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.31440004 lvth0=-2.5552838e-009            wvth0=-2.5254232e-008            pvth0=1.0487561e-015 k2=0.17889856                 lk2=-1.1186837e-008            wk2=-7.5330083e-008 pk2=3.5364757e-015             cit=0.0013910594               lcit=1.4774934e-010 wcit=-1.4808624e-009            pcit=4.7436955e-017             voff=-0.064535961 lvoff=-4.8977129e-009            wvoff=-1.6066064e-008            pvoff=4.8276534e-016 eta0=0.0042094156               weta0=1.7056591e-009             etab=-0.044952508 wetab=9.9790014e-009             u0=0.00034321299              wu0=1.1383502e-008 ua=-2.2695047e-009            lua=4.3139573e-017             wua=5.1491246e-016 pua=-2.2441249e-023            ub=1.3277369e-018             lub=-6.2097147e-027 wub=3.6121347e-025             pub=-1.4854195e-032            uc=3.0933333e-011 luc=-1.3804e-018               wuc=8.79424e-017               puc=-3.9244296e-024 vsat=107295.67                  wvsat=-0.012034691               a0=19.289417 la0=-1.2114462e-006            wa0=-7.5589616e-006            pa0=3.989891e-013 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.96776721                lketa=3.6596642e-008 wketa=3.9791849e-007             pketa=-1.795947e-014             pclm=0.4995905 wpclm=1.7164309e-007             pdiblc2=0.003                      ppdiblc2=0 wpdiblc2=0                          lpdiblc2=0                          aigbacc=0.015241794 waigbacc=-5.3557838e-009            aigc=0.0057780327               laigc=7.1223917e-012 waigc=2.4960176e-010             paigc=-1.2822495e-017            aigsd=0.0049809652 laigsd=6.0191872e-012             waigsd=8.39836e-011               paigsd=-3.6254404e-018 bigsd=0.0001728                  tvoff=0.0022887                  ltvoff=-4.98927e-013 wtvoff=-1.00771e-010              ptvoff=-1.39881e-017              kt1=-0.27731467 lkt1=4.8491675e-009             wkt1=8.4346196e-008             pkt1=-3.8364815e-015 kt2=-0.13471564                wkt2=4.3900205e-008             ute=-2.7743467 wute=8.4754488e-007             ua1=2.9346543e-009             lua1=-1.3747512e-016 wua1=-2.4855044e-015            pua1=1.1721643e-022             ub1=-6.3187283e-018 lub1=3.0570319e-025             wub1=5.7986734e-024             pub1=-2.6549974e-031 uc1=1.9577778e-010             luc1=2.0309333e-018             wuc1=2.3817733e-016 puc1=-1.0465146e-023            at=31712.018                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=5.1613245e-010 pu0=-4.4453378e-016            lvsat=-0.00013607947             pvsat=8.9769332e-010 lpclm=6.5462922e-009             ppclm=-5.411393e-015             laigbacc=-2.0387477e-010 paigbacc=2.5737717e-016             lkt2=3.5621539e-009             pkt2=-1.9236246e-015 lute=7.565187e-008              pute=-3.9538628e-014            lat=0.0011463413 leta0=4.422423e-010              peta0=-1.115163e-016             letab=1.8083096e-009 petab=-4.2886357e-016            wat=-0.021945314               pat=1.0713289e-009 vsat_ss=-1000.05                   vsat_ff=6666.71                    wvsat_ss=-6.7e-09 wvsat_ff=3.3e-08                    a0_ss=0.600003                   a0_ff=3.52333 a0_sf=-3.52333                   a0_fs=-0.600003                  la0_ss=0.0 la0_ff=-1.7969e-07                la0_sf=1.7969e-07                 la0_fs=0.0 wa0_ss=0.0                        wa0_ff=-1.92374e-06               wa0_sf=1.92374e-06 wa0_fs=0.0                        pa0_ss=5.2e-19                    pa0_ff=9.81107e-14 pa0_sf=-9.81107e-14               pa0_fs=-5.2e-19                   pdiblc2_ss=-0.00149993 pdiblc2_fs=0.00149993                 ppdiblc2_ss=7e-22                      ppdiblc2_fs=-7e-22 wpdiblc2_ss=5e-14                      wpdiblc2_fs=-5e-14                     lpdiblc2_ss=0.0 lpdiblc2_fs=0.0                        lvsat_ss=3.3e-10                    lvsat_ff=-0.000238 pvsat_ss=-2e-16                     pvsat_ff=-6e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.14 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.56101713 lvth0=7.8026342e-009             wvth0=6.9534037e-008             pvth0=-2.9323512e-015 k2=0.045062694                lk2=-5.5657305e-009            wk2=1.4483297e-008 pk2=-2.3568626e-016            cit=-0.015163493               lcit=8.4304053e-010 wcit=2.9550387e-009             pcit=-1.3887089e-016            voff=-0.22737906 lvoff=1.9416975e-009             wvoff=4.9383477e-008             pvoff=-2.2661154e-015 eta0=0.0010316576               weta0=7.0272459e-010             etab=-0.014642718 wetab=3.0366004e-010             u0=0.017862474                wu0=2.0598216e-009 ua=-1.6140415e-009            lua=1.5610118e-017             wua=1.3662389e-016 pua=-6.5531289e-024            ub=1.5608496e-018             lub=-1.6000449e-026 wub=2.0896469e-025             pub=-8.4597464e-033            uc=8.1013908e-011 luc=-3.4837841e-018            wuc=-4.0782601e-017            puc=1.4820204e-024 vsat=36128.617                  wvsat=0.024148563                a0=-31.393721 la0=9.1724559e-007             wa0=2.1872972e-005             pa0=-8.371521e-013 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.58989928                lketa=2.0726189e-008 wketa=-1.1752758e-008            pketa=-7.5327744e-016            pclm=1.6763673 wpclm=-4.3042469e-007            pdiblc2=0.017788889                lpdiblc2=-6.2113333e-010 aigbacc=0.011399206                waigbacc=2.4701738e-009             aigc=0.006100583 laigc=-6.4247222e-012            waigc=-2.4651495e-010            paigc=8.0144072e-018 aigsd=0.0050912444               laigsd=1.3874587e-012             waigsd=2.7593655e-011 paigsd=-1.2570627e-018            bigsd=0.0001728                  tvoff=0.00660097 ltvoff=-1.81614e-010              wtvoff=-2.61881e-009              ptvoff=9.17694e-017 kt1=0.24807941                 lkt1=-1.7217384e-008            wkt1=-1.8012644e-007 pkt1=7.2713693e-015             kt2=-0.080870322               wkt2=4.2313119e-009 ute=-0.60162944                wute=-4.9087432e-007            ua1=-1.7720784e-009 lua1=6.0207655e-017             wua1=1.5440785e-015             pua1=-5.2026053e-023 ub1=2.3549826e-018             lub1=-5.8592667e-026            wub1=-2.0393728e-024 pub1=6.3698203e-032             uc1=4.8553613e-010             luc1=-1.0138917e-017 wuc1=-7.0206204e-017            puc1=2.486963e-024              at=-72960.472 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=-2.1967651e-010            pu0=-5.2939184e-017            lvsat=0.0028529366 pvsat=-6.2200335e-010            lpclm=-4.2878331e-008            ppclm=1.9875454e-014 wpdiblc2=-1.0076733e-008            ppdiblc2=4.232228e-016              laigbacc=-4.2486033e-011 paigbacc=-7.1313042e-017            lkt2=1.3006506e-009             pkt2=-2.5753107e-016 lute=-1.5602253e-008            pute=1.6674978e-014             lat=0.0055425859 leta0=5.7570814e-010             peta0=-6.9393049e-017            letab=5.3529845e-010 petab=-2.2499231e-017            wat=0.04818872                 pat=-1.8743006e-009 vth0_mc=-0.0166833                 lvth0_mc=7.007e-10                  wvth0_mc=1.51151e-08 pvth0_mc=-6.34834e-16               cit_mcl=0.00722944                 cit_mc=-0.00922778 lcit_mcl=-3.03637e-10               lcit_mc=3.87567e-10                wcit_mcl=-6.54988e-09 wcit_mc=5.03837e-09                pcit_mcl=2.75095e-16                pcit_mc=-2.11611e-16 voff_ss=0.00733338                 voff_sf=0.00733338                 voff_mc=-0.0829277 voff_mcl=0.00722944                 lvoff_ss=-3.08e-10                  lvoff_sf=-3.08e-10 lvoff_mc=3.48297e-09                lvoff_mcl=-3.03637e-10               wvoff_ss=3.3e-14 wvoff_sf=3.3e-14                    wvoff_mc=3.52686e-08                wvoff_mcl=-6.54988e-09 pvoff_ss=2e-22                      pvoff_sf=2e-22                      pvoff_mc=-1.48128e-15 pvoff_mcl=2.75095e-16                eta0_mc=-0.00495611                eta0_mcl=-0.0156628 weta0_mc=5.0384e-10                 weta0_mcl=6.54987e-09                u0_ss=0.00257889 u0_ff=-0.000733338               u0_sf=-0.00138417                u0_fs=0.00184556 wu0_ss=-1.00768e-09               wu0_ff=-3.3e-15                   wu0_sf=7.55755e-10 wu0_fs=-1.00767e-09               vsat_ss=-12000                     vsat_ff=12000 vsat_sf=-5561.11                   vsat_mc=27561.1                    vsat_mcl=64594.4 wvsat_ss=-3.67e-08                  wvsat_ff=3.67e-08                   wvsat_sf=0.00503837 wvsat_mc=-0.0050384                 wvsat_mcl=-0.0352686                 a0_ss=2.8 a0_ff=-3.52333                   a0_sf=3.52333                    a0_fs=-2.8 la0_ss=-9.24e-08                  la0_ff=1.1627e-07                 la0_sf=-1.1627e-07 la0_fs=9.24e-08                   wa0_ss=0.0                        wa0_ff=1.92374e-06 wa0_sf=-1.92374e-06               wa0_fs=0.0                        pa0_ss=1.6e-19 pa0_ff=-6.34834e-14               pa0_sf=6.34834e-14                pa0_fs=-1.6e-19 pdiblc2_ss=-0.00700003                pdiblc2_fs=0.00700003                 lpdiblc2_ss=2.31e-10 lpdiblc2_fs=-2.31e-10                  lu0_ss=-1.08314e-10               lu0_ff=3.08e-11 lu0_sf=5.8135e-11                 lu0_fs=-7.75133e-11               pu0_ss=4.23223e-17 pu0_ff=-2e-23                     pu0_sf=-3.17417e-17               pu0_fs=4.23223e-17 lvsat_ss=0.000462                   lvsat_ff=-0.000462                  lvsat_sf=0.000233567 lvsat_mc=-0.00115757                lvsat_mcl=-0.00271297                pvsat_ss=-6e-16 pvsat_ff=6e-16                      pvsat_sf=-2.11611e-10               pvsat_mc=2.11608e-10 pvsat_mcl=1.48128e-09                wpdiblc2_ss=0.0                        wpdiblc2_fs=0.0 ppdiblc2_ss=1e-22                      ppdiblc2_fs=-1e-22                     leta0_mc=2.08157e-10 leta0_mcl=6.57836e-10                peta0_mc=-2.11607e-17               peta0_mcl=-2.75095e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.15 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.37656973 lvth0=-6.75461e-010              wvth0=4.1450669e-009             pvth0=1.3676593e-015 k2=0.034458006                lk2=-2.1278103e-008            wk2=-1.2222157e-009 pk2=9.1612663e-016             cit=0.0011331657               lcit=7.4814943e-011 wcit=-2.2349401e-010            pcit=-4.0848988e-017            voff=-0.11917404 lvoff=4.3968682e-012             wvoff=-1.6169444e-010            pvoff=-1.4775244e-018 eta0=0.0099656222               weta0=9.4882667e-012             etab=-0.0068677533 wetab=1.33952e-012               u0=0.010643111                wu0=1.7302133e-010 ua=5.1734187e-010             lua=-2.8484631e-016            wua=-7.6596182e-017 pua=2.1206774e-023             ub=9.9809514e-019             lub=-8.1967549e-028 wub=4.5292958e-026             pub=1.126155e-032              uc=5.3047375e-010 luc=-4.381177e-016             wuc=-4.937775e-017             puc=4.2529569e-023 vsat=101113.84                  wvsat=0.0023899269               a0=1.7142528 la0=-6.1697962e-007            wa0=6.2421997e-008             pa0=1.4861675e-013 ags=1.3309794                  lags=2.7564915e-007             wags=1.7323554e-008 pags=7.9844423e-014             keta=0.0032379996               lketa=-2.5133615e-008 wketa=-1.2223198e-008            pketa=9.5416015e-015             pclm=0.14 wpclm=6.18081e-016               pdiblc2=0.00022281481              lpdiblc2=1.5941351e-009 aigbacc=0.012372978                waigbacc=-2.5060187e-010            aigc=0.0059783326 laigc=-5.7766628e-012            waigc=2.8323628e-012             paigc=-1.6919851e-018 aigsd=0.0052776505               laigsd=5.2240303e-011             waigsd=-5.5985614e-011 paigsd=-2.8523205e-017            bigsd=0.00070743511              wbigsd=-1.4755929e-010 tvoff=0.00281494                 ltvoff=9.42842e-011               wtvoff=-5.76713e-011 ptvoff=-6.69672e-017              kt1=-0.1403084                 lkt1=5.568956e-012 wkt1=1.4512564e-009             pkt1=-9.8705525e-019            kt2=-0.078232022 wkt2=1.2563581e-009             ute=-0.85296111                wute=1.0325467e-009 ua1=8.2913889e-010             lua1=7.1726316e-017             wua1=8.873934e-017 pua1=-3.8946415e-023            ub1=-2.3548351e-019            lub1=-1.4480374e-026 wub1=-7.8573779e-026            pub1=1.6692022e-034             uc1=8.2935368e-010 luc1=-2.6409505e-016            wuc1=-2.9667887e-018            puc1=2.6692198e-023 at=90000                      jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=0 pu0=0                          lvsat=0                          pvsat=0 lpclm=2.0148096e-014             ppclm=-5.5608747e-021            lat=0 leta0=0                          peta0=0                          wat=0 pat=0                          ags_ss=-0.388711                  ags_ff=0.388711 ags_sf=0.310969                   ags_fs=-0.310969                  lags_ss=3.48675e-07 lags_ff=-3.48675e-07               lags_sf=-2.78939e-07               lags_fs=2.78939e-07 wags_ss=1.7e-13                    wags_ff=-1.7e-13                   wags_sf=2.6e-13 wags_fs=-2.6e-13                   pags_ss=-3.1e-19                   pags_ff=3.1e-19 pags_sf=-3.5e-19                   pags_fs=3.5e-19 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.16 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.37894474 lvth0=1.4549246e-009             wvth0=6.8439342e-009             pvth0=-1.0532247e-015 k2=0.0077423111               lk2=2.6858753e-009             wk2=1.8298548e-009 pk2=-1.8215806e-015            cit=0.0016233941               lcit=-3.6491997e-010 wcit=-3.461021e-010             pcit=6.9130469e-017             voff=-0.11334425 lvoff=-5.2249314e-009            wvoff=1.7977703e-010             pvoff=-3.0777743e-016 eta0=0.0099656222               weta0=9.4882667e-012             etab=-0.0068677533 wetab=1.33952e-012               u0=0.0090789864               wu0=2.38442e-010 ua=3.4013589e-010             lua=-1.2589255e-016            wua=-9.9209479e-017 pua=4.1490902e-023             ub=1.1072455e-018             lub=-9.8727521e-026 wub=6.7329951e-026             pub=-8.5056331e-033            uc=4.7675257e-011 luc=-5.0474501e-018            wuc=2.5061526e-018             puc=-4.0102914e-024 vsat=108492.55                  wvsat=-0.0016388486              a0=-0.014442242 la0=9.3365982e-007             wa0=5.7409793e-007             pa0=-3.1035657e-013 ags=0.53147285                 lags=9.9280648e-007             wags=1.8345999e-007 pags=-6.9179959e-014            keta=0.046687281                lketa=-6.4107621e-008 wketa=-1.9185867e-008            pketa=1.5787115e-014             pclm=-0.22752084 wpclm=-6.1835849e-008            pdiblc2=0.00074755015              lpdiblc2=1.1234475e-009 aigbacc=0.013384677                waigbacc=-4.3743886e-010            aigc=0.0059484398 laigc=2.103716e-011              waigc=5.4335838e-012             paigc=-4.0252803e-018 aigsd=0.0058086576               laigsd=-4.2407308e-010            waigsd=-2.1831021e-010 paigsd=1.1708196e-016             bigsd=0.001238506                wbigsd=-2.9413485e-010 tvoff=0.0028686                  ltvoff=4.61559e-011               wtvoff=-7.32303e-011 ptvoff=-5.30108e-017              kt1=-0.14672531                lkt1=5.7615379e-009 wkt1=5.7599039e-009             pkt1=-3.8658438e-015            kt2=-0.090172043 wkt2=4.6532432e-009             ute=-0.92638721                wute=7.0860794e-008 ua1=9.455976e-010              lua1=-3.2737142e-017            wua1=-2.5050022e-017 pua1=6.3122643e-023             ub1=-5.4768787e-019            lub1=2.6556693e-025 wub1=2.6510134e-025             pub1=-3.0810966e-031            uc1=6.1810844e-010 luc1=-7.4608075e-017            wuc1=3.3443349e-017             puc1=-5.9676956e-024 at=89999.997                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=1.4030199e-009 pu0=-5.868234e-017             lvsat=-0.0066187026              pvsat=3.6138116e-009 lpclm=3.2966621e-007             ppclm=5.5466751e-014             wpdiblc2=3.4567616e-010 ppdiblc2=-3.1007152e-016            laigbacc=-9.0749397e-010            paigbacc=1.6759278e-016 lbigsd=-4.7637058e-010            pbigsd=1.3147828e-016             lkt2=1.0710199e-008 pkt2=-3.0470059e-015            lute=6.5863208e-008             pute=-6.2635938e-014 lat=2.6730601e-009             leta0=0                          peta0=0 wat=0                          pat=0                          ags_ss=-0.0794664 ags_ff=0.198667                   ags_sf=0.0993333                  ags_fs=-0.0993333 lags_ss=7.12814e-08                lags_ff=-1.78204e-07               lags_sf=-8.9102e-08 lags_fs=8.9102e-08                 wags_ss=4e-15                      wags_ff=4.9e-13 wags_sf=4.4e-14                    wags_fs=-4.4e-14                   pags_ss=3.7e-20 pags_ff=7e-21                      pags_sf=4e-21                      pags_fs=-4e-21 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.17 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.3726788 lvth0=-1.3459524e-009            wvth0=3.7798467e-009             pvth0=3.1642244e-016 k2=0.021717881                lk2=-3.5612045e-009            wk2=-1.9856739e-009 pk2=-1.1603924e-016            cit=-0.0026485798              lcit=1.5446524e-009 wcit=3.0487305e-010             pcit=-2.2185543e-016            voff=-0.12535096 lvoff=1.4206924e-010             wvoff=-3.1050932e-011            pvoff=-2.1353734e-016 eta0=0.0099656222               weta0=9.4882667e-012             etab=-0.0068677533 wetab=1.33952e-012               u0=0.010959253                wu0=4.1706871e-010 ua=1.0018598e-009             lua=-4.2168312e-016            wua=3.0048282e-017 pua=-1.6287317e-023            ub=3.8588181e-019             lub=2.2372203e-025 wub=5.6146651e-026             pub=-3.5066981e-033            uc=1.4237228e-011 luc=9.899349e-018              wuc=-4.1878533e-018            puc=-1.0180708e-024 vsat=87550.122                  wvsat=0.015096282                a0=4.4289944 la0=-1.0525564e-006            wa0=-3.6017152e-007            pa0=1.0726188e-013 ags=3.4374993                  lags=-3.0618736e-007            wags=5.4814769e-008 pags=-1.1675546e-014            keta=-0.14715005                lketa=2.2537668e-008 wketa=3.1231669e-008             pketa=-6.7495232e-015            pclm=0.37663598 wpclm=1.113979e-007              pdiblc2=0.0044085574               lpdiblc2=-5.1302273e-010 aigbacc=0.012190994                waigbacc=-5.1924289e-010            aigc=0.0059611033 laigc=1.537657e-011              waigc=8.205034e-012              paigc=-5.2641185e-018 aigsd=0.004944222                laigsd=-3.7670351e-011            waigsd=-2.1232977e-011 paigsd=2.8988435e-017             bigsd=0.00029477719              wbigsd=-6.6599546e-011 tvoff=0.00445359                 ltvoff=-6.62335e-010              wtvoff=-3.52139e-010 ptvoff=7.16612e-017               kt1=-0.04826503                lkt1=-3.8250206e-008 wkt1=-1.8655835e-008            pkt1=7.0479915e-015             kt2=-0.059854191 wkt2=-5.1465618e-009            ute=-0.68660175                wute=-1.1278382e-007 ua1=3.1170134e-010             lua1=2.5061449e-016             wua1=3.5413957e-016 pua1=-1.063751e-022             ub1=9.1342042e-019             lub1=-3.8754847e-025 wub1=-1.0292726e-024            pub1=2.7047549e-031             uc1=5.850441e-010 luc1=-5.9828314e-017            wuc1=1.460592e-017              puc1=2.4526354e-024 at=55523.787                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=5.6254058e-010 pu0=-1.3852848e-016            lvsat=0.0027425645               pvsat=-3.8667915e-009 lpclm=5.9608113e-008             ppclm=-2.1968734e-014            wpdiblc2=-6.6476184e-010 ppdiblc2=1.4159427e-016             laigbacc=-3.7391792e-010            paigbacc=2.0415918e-016 lbigsd=-5.4523804e-011            pbigsd=2.9769997e-017             lkt2=-2.8418811e-009 pkt2=1.3335069e-015             lute=-4.1320891e-008            pute=1.9453202e-014 lat=0.015410869                leta0=0                          peta0=0 wat=0.024583001                pat=-1.0988602e-008            vsat_ss=-9142.99 vsat_ff=1820.51                    vsat_sf=8252.95                    vsat_fs=-6391.98 wvsat_ss=0.00101609                 wvsat_ff=-1.1e-09                   wvsat_sf=-0.00152414 wvsat_fs=0.000508048                ags_ss=-0.302308                  ags_ff=-0.0179497 ags_sf=0.173076                   ags_fs=-0.173076                  lags_ss=1.70892e-07 lags_ff=-8.13761e-08               lags_sf=-1.22065e-07               lags_fs=1.22065e-07 wags_ss=-1.78e-13                  wags_ff=-5.6e-13                   wags_sf=2.2e-13 wags_fs=-2.2e-13                   pags_ss=-6.9e-20                   pags_ff=-2.7e-20 pags_sf=-1.3e-20                   pags_fs=1.3e-20                    lvsat_ss=0.00408693 lvsat_ff=-0.000813767               lvsat_sf=-0.00368909                lvsat_fs=0.00285724 pvsat_ss=-4.54195e-10               pvsat_ff=2.7e-16                    pvsat_sf=6.81292e-10 pvsat_fs=-2.27101e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.18 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.37171248 lvth0=-1.5517795e-009            wvth0=3.2136271e-009             pvth0=4.3702721e-016 k2=0.023562007                lk2=-3.9540033e-009            wk2=-4.1597413e-009 pk2=3.4703711e-016             cit=0.0063106136               lcit=-3.6365581e-010 wcit=-1.2191846e-009            pcit=1.0276885e-016             voff=-0.097614527 lvoff=-5.765791e-009             wvoff=-4.9393462e-009            pvoff=8.3192956e-016 eta0=0.0099656219               weta0=9.4883437e-012             etab=-0.0068677423 wetab=1.3286138e-012             u0=0.011613887                wu0=1.1863577e-010 ua=-8.2746724e-010            lua=-3.2036469e-017            wua=-2.8201589e-017 pua=-3.8800946e-024            ub=1.5150141e-018             lub=-1.6783138e-026 wub=3.5945116e-026             pub=7.9622903e-034             uc=8.017987e-011 luc=-4.1464338e-018            wuc=-1.1158401e-017            puc=4.6665588e-025 vsat=100851.58                  wvsat=-0.0064371892              a0=0.12425398 la0=-1.3564664e-007            wa0=3.5541264e-007             pa0=-4.5157546e-014 ags=2.6904762                  lags=-1.4707143e-007            wags=0 pags=0                          keta=0.096098786                lketa=-2.9274335e-008 wketa=-1.922768e-008             pketa=3.9983182e-015             pclm=0.49234436 wpclm=3.4634327e-008             pdiblc2=0.0027058201               lpdiblc2=-1.5033968e-010 aigbacc=0.010978916                waigbacc=4.3925093e-010             aigc=0.0060564076 laigc=-4.9232269e-012            waigc=-1.9764821e-011            paigc=6.9346049e-019 aigsd=0.0047091174               laigsd=1.2406929e-011             waigsd=1.0872569e-010 paigsd=1.307239e-018              bigsd=6.213836e-005              wbigsd=6.0421256e-011 tvoff=0.00128854                 ltvoff=1.18201e-011               wtvoff=-3.35042e-011 ptvoff=3.79209e-018               kt1=-0.26615105                lkt1=8.1595155e-009 wkt1=2.4995884e-008             pkt1=-2.2498246e-015            kt2=-0.078290996 wkt2=2.2142877e-009             ute=-0.79470045                wute=-3.1026722e-008 ua1=2.2763185e-009             lua1=-1.6784898e-016            wua1=-2.8179988e-016 pua1=2.9079998e-023             ub1=-1.7547107e-018            lub1=1.8076346e-025 wub1=4.7390622e-025             pub1=-4.9701597e-032            uc1=2.97548e-010 luc1=1.408356e-018              wuc1=3.5762792e-017             puc1=-2.0537784e-024 at=176151.95                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=4.2310362e-010 pu0=-7.4962262e-017            lvsat=-9.0645396e-005            pvsat=7.1983775e-010 lpclm=3.4962229e-008             ppclm=-5.618093e-015             wpdiblc2=-3.8537778e-010 ppdiblc2=8.2085467e-017             laigbacc=-1.1574521e-010            paigbacc=-8.4157979e-031 lbigsd=-4.9717333e-012            pbigsd=2.7145664e-018             lkt2=1.0851584e-009 pkt2=-2.3435401e-016            lute=-1.8295867e-008            pute=2.0389414e-015 lat=-0.01028293                leta0=5.9482222e-017             peta0=-1.6417093e-023 letab=-2.3426844e-015            petab=2.3230187e-021             wat=-0.044059817 pat=3.6323186e-009             vsat_ss=19741.8                    vsat_ff=-8245.02 vsat_sf=-13209.6                   vsat_fs=13251.9                    wvsat_ss=-0.00188702 wvsat_ff=0.000770758                wvsat_sf=0.00167441                 wvsat_fs=-0.000943514 ags_ss=0.845239                   ags_ff=-0.676193                  ags_sf=-0.676193 ags_fs=0.676193                   lags_ss=-7.35362e-08               lags_ff=5.88281e-08 lags_sf=5.88281e-08                lags_fs=-5.88281e-08               wags_ss=-4.4e-13 wags_ff=-4.4e-13                   wags_sf=-4.4e-13                   wags_fs=4.4e-13 pags_ss=-3.3e-20                   pags_ff=-1.3e-20                   pags_sf=-1.3e-20 pags_fs=1.3e-20                    pdiblc2_ss=0.00103571                 pdiblc2_fs=-0.00103571 lpdiblc2_ss=-2.20607e-10               lpdiblc2_fs=2.20607e-10                lvsat_ss=-0.00206553 lvsat_ff=0.00133018                 lvsat_sf=0.000882431                lvsat_fs=-0.00132691 pvsat_ss=1.64171e-10                pvsat_ff=-1.64171e-10               pvsat_sf=-6e-16 pvsat_fs=8.20857e-11                wpdiblc2_ss=-3.3e-16                   wpdiblc2_fs=3.3e-16 ppdiblc2_ss=-2e-22                     ppdiblc2_fs=2e-22 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.19 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.40441375 lvth0=1.2932317e-009             wvth0=1.5294168e-008             pvth0=-6.1397987e-016 k2=0.019198258                lk2=-3.5743571e-009            wk2=-2.8468381e-012 pk2=-1.4612709e-017            cit=-0.00021967391             lcit=2.044792e-010 wcit=3.0302341e-010             pcit=-2.9663243e-017            voff=-0.15827866 lvoff=-4.8801164e-010            wvoff=1.4893003e-008             pvoff=-8.9348486e-016 eta0=0.0041872917               weta0=1.6043075e-009             etab=-0.0055377484 wetab=-9.1444169e-010            u0=0.015951324                wu0=-6.3536129e-010 ua=-1.2455457e-009            lua=4.33636e-018               wua=-7.8508693e-017 pua=4.9662342e-025             ub=1.2964798e-018             lub=2.229346e-027 wub=1.1369734e-025             pub=-5.9682146e-033            uc=1.273598e-011 luc=1.7211846e-018             wuc=3.3884414e-018             puc=-7.9891941e-025 vsat=80535.239                  wvsat=0.003349474                a0=0.33660924 la0=-1.5412155e-007            wa0=6.0612962e-007             pa0=-6.6969924e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.33606625                lketa=8.3240227e-009 wketa=5.9573104e-008             pketa=-2.8573501e-015            pclm=1.3271838 wpclm=-1.9565526e-007            pdiblc2=-0.0033351852              lpdiblc2=3.7522778e-010 aigbacc=0.009817787                waigbacc=1.7278878e-010             aigc=0.0060314114 laigc=-2.7485605e-012            waigc=2.0354712e-011             paigc=-2.7969388e-018 aigsd=0.0048614584               laigsd=-8.4674106e-013            waigsd=8.4224138e-011 paigsd=3.4388741e-018             bigsd=7.7558704e-005             wbigsd=5.2001748e-011 tvoff=0.00108567                 ltvoff=2.94702e-011               wtvoff=7.96676e-011 ptvoff=-6.05386e-018              kt1=-0.17129118                lkt1=-9.3293233e-011 wkt1=-7.9614067e-009            pkt1=6.1745968e-016             kt2=-0.093596509 wkt2=4.5169266e-009             ute=-0.5593113                 wute=-1.4287748e-007 ua1=1.5165462e-009             lua1=-1.0174879e-016            wua1=-1.6317655e-016 pua1=1.8759768e-023             ub1=-1.2281461e-018            lub1=1.3495234e-025 wub1=2.7272292e-025             pub1=-3.2198649e-032            uc1=3.8281619e-010 luc1=-6.0099768e-018            wuc1=5.3783588e-018             puc1=5.8966731e-025 at=68103.302                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=4.5746623e-011 pu0=-9.3645181e-018            lvsat=0.0016768761               pvsat=-1.3160195e-010 lpclm=-3.7668801e-008            ppclm=1.4417101e-014             wpdiblc2=2.1395111e-009 ppdiblc2=-1.3757987e-016            laigbacc=-1.4727006e-011            paigbacc=2.3182207e-017 lbigsd=-6.3133032e-012            pbigsd=3.4470636e-018             lkt2=2.416738e-009 pkt2=-4.3468359e-016            lute=-3.8774724e-008            pute=1.1769958e-014 lat=-0.00088269765             leta0=5.0271479e-010             peta0=-1.3874928e-016 letab=-1.1571181e-010            petab=7.9674339e-017             wat=-0.0068751903 pat=3.9725611e-010             vsat_ss=-5353.72                   vsat_ff=11294.5 vsat_sf=-7411.11                   vsat_fs=-4833.33                   wvsat_ss=-0.00158138 wvsat_ff=-0.00111626                wvsat_sf=0.00404647                 wvsat_fs=-4.4e-09 a0_ss=-0.850001                  a0_sf=0.868889                   a0_fs=0.850001 la0_ss=7.39497e-08                la0_sf=-7.55933e-08               la0_fs=-7.39497e-08 wa0_ss=-3.3e-13                   wa0_sf=-4.74413e-07               wa0_fs=3.3e-13 pa0_ss=-4e-20                     pa0_sf=4.1274e-14                 pa0_fs=4e-20 pdiblc2_ss=-0.0015                    pdiblc2_fs=0.0015                     lpdiblc2_ss=-3.3e-16 lpdiblc2_fs=3.3e-16                    lvsat_ss=0.000117772                lvsat_ff=-0.000369749 lvsat_sf=0.000377967                lvsat_fs=0.0002465                  pvsat_ss=1.3758e-10 pvsat_ff=2e-16                      pvsat_sf=-2.0637e-10                pvsat_fs=-1.3e-16 wpdiblc2_ss=6.7e-15                    wpdiblc2_fs=-6.7e-15                   ppdiblc2_ss=-1e-22 ppdiblc2_fs=1e-22 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.20 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.35997891 lvth0=-9.7294525e-010            wvth0=-3.681667e-010             pvth0=1.8479921e-016 k2=0.073868782                lk2=-6.3625538e-009            wk2=-1.7983824e-008 pk2=9.0241711e-016             cit=0.0011902688               lcit=1.3257212e-010 wcit=-1.3712307e-009            pcit=5.5723715e-017             voff=-0.075423109 lvoff=-4.7136446e-009            wvoff=-1.0121681e-008            pvoff=3.8226405e-016 eta0=0.0093777778               weta0=-1.1162667e-009            etab=-0.032908866 wetab=3.4031731e-009             u0=0.026337765                wu0=-2.8095233e-009 ua=-8.9077829e-010            lua=-1.3756779e-017            wua=-2.3787214e-016 pua=8.6241594e-024             ub=2.0834535e-018             lub=-3.7906313e-026 wub=-5.1407801e-026            pub=2.4521476e-033             uc=3.0522621e-010 luc=-1.3195817e-017            wuc=-6.1821508e-017            puc=2.526788e-024 vsat=99571.52                   wvsat=-0.0078173072              a0=10.304307 la0=-6.6247414e-007            wa0=-2.6530916e-006            pa0=9.9250359e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.3779993                 lketa=1.0462609e-008 wketa=7.5905212e-008             pketa=-3.6902876e-015            pclm=0.87247107 wpclm=-3.1949699e-008            pdiblc2=0.0040222222               ppdiblc2=0 lpdiblc2=0                          aigbacc=-0.0053667704              waigbacc=5.8964926e-009 aigc=0.006418962                laigc=-2.2513642e-011            waigc=-1.0034565e-010 paigc=3.3587794e-018             aigsd=0.0041095766               laigsd=3.749923e-011 waigsd=5.5976174e-010             paigsd=-2.0813544e-017            bigsd=-0.0010683788 wbigsd=6.7768363e-010             tvoff=0.00292794                 ltvoff=-6.44856e-011 wtvoff=-4.49791e-010              ptvoff=2.09486e-017               kt1=-0.10099019 lkt1=-3.6786434e-009            wkt1=-1.1926967e-008            pkt1=8.1970328e-016 kt2=-0.013897074               wkt2=-2.2066732e-008            ute=-2.0628444 wute=4.5906467e-007             ua1=-4.7913018e-009            lua1=2.1995146e-016 wua1=1.7328677e-015             pua1=-7.7938487e-023            ub1=9.3803975e-018 lub1=-4.0608339e-025            wub1=-2.7730493e-024            pub1=1.2313573e-031 uc1=5.3250916e-010             luc1=-1.3644318e-017            wuc1=5.4322001e-017 puc1=-1.9064584e-024            at=-23253.577                 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-4.8396191e-010 pu0=1.0151774e-016             lvsat=0.00070602572              pvsat=4.3790389e-010 lpclm=-1.4478452e-008            ppclm=6.0681175e-015             wpdiblc2=-5.5813333e-010 laigbacc=7.5968542e-010             paigbacc=-2.6872669e-016            lbigsd=5.212951e-011 pbigsd=-2.8462713e-017            lkt2=-1.6479332e-009            pkt2=9.2108297e-016 lute=3.7905467e-008             pute=-1.8929092e-014            lat=0.0037765032 leta0=2.38e-010                  peta0=2.9385381e-030             letab=1.2802152e-009 petab=-1.4052402e-016            wat=0.0080659009               pat=-3.6473955e-010 u0_ss=0.00190815                 u0_ff=-0.000954074               wu0_ss=-1.04185e-09 wu0_ff=5.20924e-10                vsat_ss=1725.95                    vsat_ff=3940.72 vsat_sf=-9540.74                   vsat_fs=9540.74                    wvsat_ss=-0.00148834 wvsat_ff=0.00148835                 wvsat_sf=0.00520924                 wvsat_fs=-0.00520924 a0_ss=3.46222                    a0_ff=-2.86222                   a0_sf=-0.613336 a0_fs=-3.46222                   la0_ss=-1.45974e-07               la0_ff=1.45973e-07 la0_sf=3.3e-13                    la0_fs=1.45974e-07                wa0_ss=-1.56278e-06 wa0_ff=1.56277e-06                wa0_sf=3.34883e-07                wa0_fs=1.56278e-06 pa0_ss=7.97016e-14                pa0_ff=-7.97014e-14               pa0_sf=-4e-20 pa0_fs=-7.97016e-14               pdiblc2_ss=-0.00149991                pdiblc2_fs=0.00149991 ppdiblc2_ss=6e-22                      ppdiblc2_fs=-6e-22                     lpdiblc2_ss=-3.3e-16 lpdiblc2_fs=3.3e-16                    lu0_ss=-9.73156e-11               lu0_ff=4.86578e-11 pu0_ss=5.31343e-17                pu0_ff=-2.65671e-17               lvsat_ss=-0.000243289 lvsat_ff=5.28922e-06                lvsat_sf=0.000486578                lvsat_fs=-0.000486578 pvsat_ss=1.32835e-10                pvsat_ff=-1.32836e-10               pvsat_sf=-2.65671e-10 pvsat_fs=2.65671e-10                wpdiblc2_ss=6.7e-15                    wpdiblc2_fs=-6.7e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.21 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.4262675 lvth0=1.8111756e-009             wvth0=-4.0392613e-009            pvth0=3.3898519e-016 k2=0.089029598                lk2=-6.9993081e-009            wk2=-9.5226331e-009 pk2=5.4704711e-016             cit=-0.010298272               lcit=6.1509083e-010 wcit=2.9862814e-010             pcit=-1.4410355e-017            voff=-0.10043056 lvoff=-3.6633315e-009            wvoff=-1.9930405e-008            pvoff=7.9423046e-016 eta0=0.0014640666               weta0=4.6662925e-010             etab=-0.017132505 wetab=1.6630837e-009             u0=0.024909091                wu0=-1.7876312e-009 ua=-1.3089513e-009            lua=3.8064892e-018             wua=-2.9955314e-017 pua=-1.0834747e-025            ub=2.0487317e-018             lub=-3.6447996e-026 wub=-5.7418918e-026            pub=2.7046146e-033             uc=1.5471944e-011 luc=-1.0261379e-018            wuc=-4.9966887e-018            puc=1.4014561e-025 vsat=45883.238                  wvsat=0.01882254                 a0=11.145195 la0=-6.9779144e-007            wa0=-1.3532765e-006            pa0=4.4658124e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.6709001                 lketa=2.2764442e-008 wketa=3.2473687e-008             pketa=-1.8661635e-015            pclm=0.73893137 wpclm=8.1415299e-008             pdiblc2=0.00035555556              lpdiblc2=1.54e-010 aigbacc=0.01894877                 waigbacc=-1.6518886e-009            aigc=0.005519132 laigc=1.5279217e-011             waigc=7.0957288e-011             paigc=-3.8359438e-018 aigsd=0.0050463575               laigsd=-1.8455688e-012            waigsd=5.2101886e-011 paigsd=5.0817029e-019             bigsd=0.0001728                  tvoff=0.00164043 ltvoff=-1.04101e-011              wtvoff=8.9651e-011                ptvoff=-1.70803e-018 kt1=-0.14669239                lkt1=-1.7591511e-009            wkt1=3.5418961e-008 pkt1=-1.1688257e-015            kt2=-0.068133585               wkt2=-2.7229465e-009 ute=-2.0081319                 wute=2.7707599e-007             ua1=2.1595468e-009 lua1=-7.1984178e-017            wua1=-6.0258888e-016            pua1=2.0150688e-023 ub1=-3.6944152e-018            lub1=1.4305875e-025             wub1=1.2635984e-024 pub1=-4.6403471e-032            uc1=2.1027467e-010             luc1=-1.1046933e-019 wuc1=8.0086552e-017             puc1=-2.9885696e-024            at=6427.7055 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=-4.2395757e-010            pu0=5.8598277e-017             lvsat=0.0029609336 pvsat=-6.8096969e-010            lpclm=-8.8697849e-009            ppclm=1.3067876e-015 wpdiblc2=-5.5813333e-010            ppdiblc2=2.050537e-031              laigbacc=-2.6156729e-010 paigbacc=4.8305324e-017             lkt2=6.3000031e-010             pkt2=1.08644e-016 lute=3.5607538e-008             pute=-1.1285568e-014            lat=0.0025298893 leta0=5.7037587e-010             peta0=-6.6481629e-017            letab=6.1760803e-010 petab=-6.7440262e-017            wat=0.0048427749               pat=-2.2936826e-010 vth0_mc=0.0222444                  lvth0_mc=-9.34267e-10               wvth0_mc=-6.13947e-09 pvth0_mc=2.57858e-16                cit_mcl=-0.00589111                lcit_mcl=2.47427e-10 wcit_mcl=6.13946e-10                pcit_mcl=-2.57858e-17               voff_ss=0.0148296 voff_ff=0.0074963                  voff_sf=0.0148296                  voff_mc=-0.0370741 voff_mcl=-0.00963926                lvoff_ss=-6.22844e-10               lvoff_ff=-3.14844e-10 lvoff_sf=-6.22844e-10               lvoff_mc=1.55711e-09                lvoff_mcl=4.04849e-10 wvoff_ss=-4.09298e-09               wvoff_ff=-4.09298e-09               wvoff_sf=-4.09298e-09 wvoff_mc=1.02324e-08                wvoff_mcl=2.66044e-09                pvoff_ss=1.71905e-16 pvoff_ff=1.71905e-16                pvoff_sf=1.71905e-16                pvoff_mc=-4.29763e-16 pvoff_mcl=-1.11738e-16               eta0_mc=-0.00628223                eta0_mcl=-0.00741481 weta0_mc=1.2279e-09                 weta0_mcl=2.04649e-09                u0_ss=-0.000425188 u0_ff=-0.000903696               u0_sf=-0.00074963                u0_fs=0.00074963 wu0_ss=6.32551e-10                wu0_ff=9.30226e-11                wu0_sf=4.09298e-10 wu0_fs=-4.09298e-10               vsat_ss=-26311                     vsat_ff=26311 vsat_sf=13207.4                    vsat_fs=-5792.59                   vsat_mc=32576.3 wvsat_ss=0.00781386                 wvsat_ff=-0.00781386                wvsat_sf=-0.00520925 wvsat_fs=0.00316275                 wvsat_mc=-0.00777665                a0_ss=-0.0622244 a0_ff=2.86222                    a0_sf=-2.86222                   a0_fs=0.0622244 la0_ss=2.05367e-09                la0_ff=-9.44533e-08               la0_sf=9.44533e-08 la0_fs=-2.05367e-09               wa0_ss=1.56278e-06                wa0_ff=-1.56277e-06 wa0_sf=1.56277e-06                wa0_fs=-1.56278e-06               pa0_ss=-5.15715e-14 pa0_ff=5.15715e-14                pa0_sf=-5.15715e-14               pa0_fs=5.15715e-14 pdiblc2_ss=-0.00700004                pdiblc2_fs=0.00700004                 lpdiblc2_ss=2.31e-10 lpdiblc2_fs=-2.31e-10                  at_mc=11244.4                    lu0_ss=6.84489e-13 lu0_ff=4.65422e-11                lu0_sf=3.14844e-11                lu0_fs=-3.14844e-11 pu0_ss=-1.71905e-17               pu0_ff=-8.59529e-18               pu0_sf=-1.71905e-17 pu0_fs=1.71905e-17                lvsat_ss=0.000934266                lvsat_ff=-0.000934266 lvsat_sf=-0.000468844               lvsat_fs=0.000157422                lvsat_mc=-0.0013682 pvsat_ss=-2.57858e-10               pvsat_ff=2.57858e-10                pvsat_sf=1.71905e-10 pvsat_fs=-8.59526e-11               pvsat_mc=3.2662e-10                 wpdiblc2_ss=-3.3e-15 wpdiblc2_fs=3.3e-15                    ppdiblc2_ss=-2e-22                     ppdiblc2_fs=2e-22 lat_mc=-0.000472267               leta0_mc=2.63853e-10                leta0_mcl=3.11422e-10 peta0_mc=-5.15715e-17               peta0_mcl=-8.59525e-17               wat_mc=-0.00613947 pat_mc=2.57858e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_mac.22 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.36655807 lvth0=-3.6900702e-009            wvth0=1.3818477e-009             pvth0=2.1996915e-015 k2=0.036083654                lk2=-2.8077385e-008            wk2=-1.6708948e-009 pk2=2.7927287e-015             cit=0.00023111811              lcit=-1.2469172e-010 wcit=2.5471122e-011             pcit=1.421485e-017              voff=-0.1234315 lvoff=-5.8275177e-009            wvoff=1.0133624e-009             pvoff=1.6081309e-015 eta0=0.010567185                weta0=-1.5654311e-010            etab=-0.0078955852 wetab=2.8502111e-010             u0=0.011413556                wu0=-3.9621333e-011 ua=3.9795887e-010             lua=-3.086736e-016             wua=-4.3646473e-017 pua=2.7783107e-023             ub=1.4169172e-018             lub=-4.8255908e-026 wub=-7.0301945e-026            pub=2.435395e-032              uc=4.5023847e-010 luc=-3.6135906e-016            wuc=-2.7232811e-017            puc=2.1344185e-023 vsat=109613.26                  wvsat=4.4088444e-005             a0=2.1211719 la0=-4.7894519e-007            wa0=-4.9887669e-008            pa0=1.1051925e-013 ags=1.4232152                  lags=4.9466262e-007             wags=-8.133534e-009 pags=1.9396705e-014             keta=-0.08853915                lketa=6.8992317e-008 wketa=1.3107295e-008             pketa=-1.6437156e-014            pclm=0.074801852 wpclm=1.7994689e-008             pdiblc2=0.00014488615              lpdiblc2=2.2952594e-009 aigbacc=0.011623333                waigbacc=-4.37e-011                 aigc=0.0059916363 laigc=-2.6091067e-011            waigc=-8.3945942e-013            paigc=3.9147906e-018 aigsd=0.0050437597               laigsd=-1.0808354e-010            waigsd=8.5682537e-012 paigsd=1.5726175e-017             bigsd=0.0001728                  tvoff=0.00247841 ltvoff=-1.93342e-010              wtvoff=3.52113e-011               ptvoff=1.24176e-017 kt1=-0.13562712                lkt1=7.376565e-013              wkt1=1.5922372e-010 pkt1=3.4638342e-019             kt2=-0.071096704               wkt2=-7.1298978e-010 ute=-0.78492963                wute=-1.7744142e-008            ua1=1.4842296e-009 lua1=-6.9835373e-017            wua1=-9.2065696e-017            pua1=1.2461095e-025 ub1=-7.0678485e-019            lub1=-3.9802279e-027            wub1=5.1505393e-026 pub1=-2.7311203e-033            uc1=9.0769646e-010             luc1=-2.8517306e-016 wuc1=-2.4589396e-017            puc1=3.2509729e-023             at=108296.3 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=0                          pu0=0                          lvsat=0 pvsat=0                          lpclm=0                          ppclm=0 wpdiblc2=2.1508313e-011             ppdiblc2=-1.9351029e-016            lat=-7.0112424e-009 leta0=0                          peta0=0                          wat=-0.005049778 pat=1.9351029e-015             ags_ss=-0.505942                  ags_ff=0.505942 ags_sf=0.404753                   ags_fs=-0.404753                  lags_ss=4.5383e-07 lags_ff=-4.5383e-07                lags_sf=-3.63064e-07               lags_fs=3.63064e-07 wags_ss=3.23556e-08                wags_ff=-3.23556e-08               wags_sf=-2.58845e-08 wags_fs=2.58845e-08                pags_ss=-2.9023e-14                pags_ff=2.9023e-14 pags_sf=2.32184e-14                pags_fs=-2.32184e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_mac.23 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.37029672 lvth0=-3.3650152e-010            wvth0=4.4570791e-009             pvth0=-5.5879105e-016 k2=0.0080761272               lk2=-2.9546335e-009            wk2=1.7377216e-009 pk2=-2.6480016e-016            cit=0.00019465172              lcit=-9.1981363e-011 wcit=4.8230807e-011             pcit=-6.200587e-018             voff=-0.1248711 lvoff=-4.5361908e-009            wvoff=3.3611893e-009             pvoff=-4.9786984e-016 eta0=0.010567185                weta0=-1.5654311e-010            etab=-0.0078955852 wetab=2.8502111e-010             u0=0.010393329                wu0=-1.2431647e-010 ua=1.077583e-010              lua=-4.8363693e-017            wua=-3.5073262e-017 pua=2.0092937e-023             ub=1.6239722e-018             lub=-2.339842e-025 wub=-7.5286627e-026            pub=2.882521e-032              uc=9.9571279e-011 luc=-4.6810594e-017            wuc=-1.1817149e-017            puc=7.5163362e-024 vsat=97315.41                   wvsat=0.0014460433               a0=1.692364 la0=-9.4304527e-008            wa0=1.0301942e-007             pa0=-2.6638408e-014 ags=1.1519585                  lags=7.3797986e-007             wags=1.2205949e-008 pags=1.1521888e-015             keta=0.0065370473               lketa=-1.6291032e-008 wketa=-8.1044022e-009            pketa=2.5897367e-015             pclm=-0.62397923 wpclm=4.7586666e-008             pdiblc2=0.003402716                lpdiblc2=-6.2701407e-010 aigbacc=0.012193654                waigbacc=-1.0871654e-010            aigc=0.005934217 laigc=2.5414068e-011             waigc=9.3590884e-012             paigc=-5.2333069e-018 aigsd=0.0049355964               laigsd=-1.1061049e-011            waigsd=2.2654694e-011 paigsd=3.0906379e-018             bigsd=0.0001728                  tvoff=0.00257692 ltvoff=-2.81707e-010              wtvoff=7.27163e-012               ptvoff=3.74795e-017 kt1=-0.11623884                lkt1=-1.739055e-008             wkt1=-2.6543618e-009 pkt1=2.5241326e-015             kt2=-0.066994347               wkt2=-1.7438009e-009 ute=-0.47454166                wute=-5.3848577e-008            ua1=1.310304e-009 lua1=8.6175917e-017             wua1=-1.2570898e-016            pua1=3.0302639e-023 ub1=4.9968824e-019             lub1=-1.0861866e-024            wub1=-2.3974469e-026 pub1=6.4974315e-032             uc1=7.6416296e-010             luc1=-1.5642351e-016 wuc1=-6.8676978e-018            puc1=1.6613365e-023             at=104102.2 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=9.1514354e-010             pu0=7.5971533e-017             lvsat=0.011031171 pvsat=-1.2575535e-009            lpclm=6.2680663e-007             ppclm=-2.6544004e-014 wpdiblc2=-3.8714963e-010            ppdiblc2=1.7305588e-016             laigbacc=-5.1157748e-010 paigbacc=5.8319833e-017             lkt2=-3.6798136e-009            pkt2=9.2463759e-016 lute=-2.7841801e-007            pute=3.2385678e-014             lat=0.0037620971 leta0=0                          peta0=0                          wat=-0.0038922083 pat=-1.0383381e-009            ags_ss=-0.135388                  ags_ff=0.338469 ags_sf=0.169235                   ags_fs=-0.169235                  lags_ss=1.21443e-07 lags_ff=-3.03607e-07               lags_sf=-1.51803e-07               lags_fs=1.51803e-07 wags_ss=1.54342e-08                wags_ff=-3.85855e-08               wags_sf=-1.92927e-08 wags_fs=1.92927e-08                pags_ss=-1.38445e-14               pags_ff=3.46112e-14 pags_sf=1.73056e-14                pags_fs=-1.73056e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_mac.24 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.37336188 lvth0=1.0336251e-009             wvth0=3.9683764e-009             pvth0=-3.4034095e-016 k2=0.015507636                lk2=-6.2765179e-009            wk2=-2.7164629e-010 pk2=6.3338726e-016             cit=-0.0023370065              lcit=1.0396699e-009 wcit=2.1887884e-010             pcit=-8.2480257e-017            voff=-0.1394312 lvoff=1.9721737e-009             wvoff=3.855096e-009              pvoff=-7.1864616e-016 eta0=0.010567185                weta0=-1.5654311e-010            etab=-0.0078955852 wetab=2.8502111e-010             u0=0.012453609                wu0=4.6264729e-012 ua=1.1475367e-009             lua=-5.1314464e-016            wua=-1.015855e-017 pua=8.9560611e-024             ub=6.4230133e-019             lub=2.0482268e-025 wub=-1.4625137e-026            pub=1.7095236e-033             uc=-7.6171348e-012 luc=1.1026272e-018             wuc=1.8439508e-018             puc=1.4098245e-024 vsat=151358.28                  wvsat=-0.0025147703              a0=2.834408 la0=-6.0479819e-007            wa0=7.9934322e-008             pa0=-1.6319371e-014 ags=3.0943679                  lags=-1.3027713e-007            wags=1.4951906e-007 pags=-6.022677e-014             keta=-0.023816795               lketa=-2.7228649e-009 wketa=-2.8083106e-009            pketa=2.2238377e-016             pclm=0.86913034 wpclm=-2.4530543e-008            pdiblc2=0.002                      lpdiblc2=0 aigbacc=0.0094391439               waigbacc=2.4026783e-010             aigc=0.005986487 laigc=2.049388e-012              waigc=1.1991541e-012             paigc=-1.5858162e-018 aigsd=0.0046631896               laigsd=1.1070478e-010             waigsd=5.6331964e-011 paigsd=-1.1963102e-017            bigsd=-3.0495318e-005            wbigsd=2.3175666e-011 tvoff=0.00306283                 ltvoff=-4.98908e-010              wtvoff=3.17102e-011 ptvoff=2.65555e-017               kt1=-0.11977538                lkt1=-1.5809718e-008 wkt1=1.0810202e-009             pkt1=8.5441684e-016             kt2=-0.080801273 wkt2=6.3483276e-010             ute=-1.2842486                 wute=5.2166703e-008 ua1=2.1475694e-009             lua1=-2.8808172e-016            wua1=-1.5256001e-016 pua1=4.2305049e-023             ub1=-4.3835778e-018            lub1=1.0966333e-024 wub1=4.3269891e-025             pub1=-1.3915868e-031            uc1=4.0981254e-010 luc1=1.9711299e-018             wuc1=6.2969832e-017             puc1=-1.4604011e-023 at=191436.07                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-5.8018732e-012 pu0=1.833404e-017              lvsat=-0.013125992               pvsat=5.1293017e-010 lpclm=-4.0613345e-008            ppclm=5.6923889e-015             laigbacc=7.1968847e-010 paigbacc=-9.7676178e-017            lbigsd=9.0873007e-011             pbigsd=-1.0359523e-017 lkt2=2.4918819e-009             pkt2=-1.3861166e-016            lute=8.3520971e-008 pute=-1.5003152e-014            lat=-0.035276144               leta0=0 peta0=0                          wat=-0.012928789               pat=3.0010137e-009 vsat_ss=-9304.84                   vsat_ff=6304.36                    vsat_sf=4652.42 vsat_fs=-7754.04                   wvsat_ss=0.00106075                 wvsat_ff=-0.00123754 wvsat_sf=-0.000530376               wvsat_fs=0.00088396                 ags_ss=-0.515043 ags_ff=-0.0305792                 ags_sf=0.294872                   ags_fs=-0.294872 lags_ss=2.91148e-07                lags_ff=-1.38642e-07               lags_sf=-2.07963e-07 lags_fs=2.07963e-07                wags_ss=5.87149e-08                wags_ff=3.48605e-09 wags_sf=-3.36154e-08               wags_fs=3.36154e-08                pags_ss=-3.31909e-14 pags_ff=1.58052e-14                pags_sf=2.37078e-14                pags_fs=-2.37078e-14 lvsat_ss=0.00415927                 lvsat_ff=-0.00281805                lvsat_sf=-0.00207963 lvsat_fs=0.00346605                 pvsat_ss=-4.74156e-10               pvsat_ff=5.53182e-10 pvsat_sf=2.37078e-10                pvsat_fs=-3.9513e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_mac.25 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.36066254 lvth0=-1.6713344e-009            wvth0=1.6384442e-010             pvth0=4.7002436e-016 k2=-0.0028058244              lk2=-2.3757509e-009            wk2=3.1177801e-009 pk2=-8.8560554e-017            cit=0.0034717531               lcit=-1.9759593e-010 wcit=-4.3565912e-010            pcit=5.6936328e-017             voff=-0.10906016 lvoff=-4.4968587e-009            wvoff=-1.7803519e-009            pvoff=4.8170426e-016 eta0=0.010567168                weta0=-1.565384e-010             etab=-0.0078956427 wetab=2.8502912e-010             u0=0.011613585                wu0=1.1871917e-010 ua=-1.0905588e-009            lua=-3.64303e-017              wua=4.4411677e-017 pua=-2.6673974e-024            ub=1.6030098e-018             lub=1.9176807e-028 wub=1.1658283e-026             pub=-3.888845e-033             uc=-1.9626766e-011 luc=3.6606787e-018             wuc=1.6388231e-017             puc=-1.6881072e-024 vsat=90331.976                  wvsat=-0.0035337792              a0=2.8246856 la0=-6.0272733e-007            wa0=-3.8990649e-007            pa0=8.3756723e-014 ags=3.5551226                  lags=-2.2841789e-007            wags=-2.3864242e-007 pags=2.2451624e-014             keta=0.080780715                lketa=-2.5002134e-008 wketa=-1.4999893e-008            pketa=2.8191908e-015             pclm=0.63620466 wpclm=-5.0711166e-009            pdiblc2=0.0010588042               lpdiblc2=2.004747e-010 aigbacc=0.014071254                waigbacc=-4.1423438e-010            aigc=0.0060133681 laigc=-3.6762926e-012            waigc=-7.8859296e-012            paigc=3.4930662e-019 aigsd=0.005125132                laigsd=1.2311039e-011             waigsd=-6.0943557e-012 paigsd=1.3337043e-018             bigsd=0.00043699988              wbigsd=-4.3040523e-011 tvoff=0.000228294                ltvoff=1.04849e-010               wtvoff=2.59124e-010 ptvoff=-2.18838e-017              kt1=-0.21868352                lkt1=5.2577173e-009 wkt1=1.1894847e-008             pkt1=-1.4489283e-015            kt2=-0.068676554 wkt2=-4.392983e-010             ute=-0.77648871                wute=-3.6053162e-008 ua1=9.9237532e-010             lua1=-4.2025386e-017            wua1=7.2568449e-017 pua1=-5.647313e-024             ub1=1.4575862e-018             lub1=-1.475346e-025 wub1=-4.1268772e-025            pub1=4.0908667e-032             uc1=4.5760342e-010 luc1=-8.2083288e-018            wuc1=-8.4125043e-018            puc1=6.0042662e-025 at=8490.5732                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=1.7312334e-010 pu0=-5.9677036e-018            lvsat=-0.00012738931             pvsat=7.2997907e-010 lpclm=8.9998235e-009             ppclm=1.547531e-015              wpdiblc2=6.9198603e-011 ppdiblc2=-1.4739303e-017            laigbacc=-2.6695098e-010            paigbacc=4.1732792e-017 lbigsd=-8.7034693e-012            pbigsd=3.7445255e-018             lkt2=-9.0683153e-011 pkt2=9.0178252e-017             lute=-2.4631874e-008            pute=3.7876794e-015 lat=0.0036912478               leta0=3.6326643e-015             peta0=-1.0026153e-021 letab=1.2252684e-014             petab=-1.705303e-021             wat=0.0022147232 pat=-2.2455448e-010            u0_ss=-0.000194356               u0_ff=0.000194356 wu0_ss=5.36423e-11                wu0_ff=-5.36423e-11               vsat_ss=21985.9 vsat_ff=-13779.5                   vsat_sf=-10711.6                   vsat_fs=15781.3 wvsat_ss=-0.00250639                wvsat_ff=0.0022983                  wvsat_sf=0.000984984 wvsat_fs=-0.00164164                ags_ss=1.44004                    ags_ff=-1.15203 ags_sf=-1.15203                   ags_fs=1.15203                    lags_ss=-1.25283e-07 lags_ff=1.00226e-07                lags_sf=1.00226e-07                lags_fs=-1.00226e-07 wags_ss=-1.64164e-07               wags_ff=1.31331e-07                wags_sf=1.31331e-07 wags_fs=-1.31331e-07               pags_ss=1.42823e-14                pags_ff=-1.14258e-14 pags_sf=-1.14258e-14               pags_fs=1.14258e-14                pdiblc2_ss=0.00176455 pdiblc2_fs=-0.00176455                lpdiblc2_ss=-3.75849e-10               lpdiblc2_fs=3.75849e-10 lu0_ss=4.13979e-11                lu0_ff=-4.13979e-11               pu0_ss=-1.14258e-17 pu0_ff=1.14258e-17                lvsat_ss=-0.00250566                lvsat_ff=0.00145982 lvsat_sf=0.00119291                 lvsat_fs=-0.00154697                pvsat_ss=2.85645e-10 pvsat_ff=-1.99952e-10               pvsat_sf=-8.56936e-11               pvsat_fs=1.42823e-10 wpdiblc2_ss=-2.01159e-10               wpdiblc2_fs=2.01159e-10                ppdiblc2_ss=4.28468e-17 ppdiblc2_fs=-4.28468e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_mac.26 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.37673715 lvth0=-2.7284304e-010            wvth0=7.6554261e-009             pvth0=-1.8174325e-016 k2=0.025694                   lk2=-4.8552356e-009            wk2=-1.7956717e-009 pk2=3.3890975e-016             cit=-0.00017842273             lcit=1.1996936e-010 wcit=2.9163808e-010             pcit=-6.3385289e-018            voff=-0.11302552 lvoff=-4.1518725e-009            wvoff=2.4031369e-009             pvoff=1.1774073e-016 eta0=0.010373844                weta0=-1.0318085e-010            etab=-0.010510707 wetab=4.5809487e-010             u0=0.014683833                wu0=-2.8553386e-010 ua=-1.4233608e-009            lua=-7.4765247e-018            wua=-2.9431736e-017 pua=3.7569796e-024             ub=1.7978146e-018             lub=-1.6756248e-026 wub=-2.4671078e-026            pub=-7.2819058e-034            uc=2.150353e-011 luc=8.2342869e-020             wuc=9.6859755e-019             puc=-3.4659909e-025 vsat=78545.957                  wvsat=0.0038985156               a0=0.92285094 la0=-4.3726771e-007            wa0=4.4432692e-007             pa0=1.1178416e-014 ags=0.82993827                 lags=8.6731481e-009             wags=4.6937037e-008 pags=-2.3937889e-015            keta=-0.29917229                lketa=8.0537772e-009 wketa=4.9390373e-008             pketa=-2.7827623e-015            pclm=0.38336074 wpclm=6.48399e-008               pdiblc2=0.0062910988               lpdiblc2=-2.5473493e-010 aigbacc=0.0093104599               waigbacc=3.1281107e-010             aigc=0.0061152847 laigc=-1.2543035e-011            waigc=-2.7943141e-012            paigc=-9.3663932e-020 aigsd=0.0049446529               laigsd=2.8012724e-011             waigsd=6.1262457e-011 paigsd=-4.5263383e-018            bigsd=5.2362161e-005             wbigsd=5.8955994e-011 tvoff=0.00125718                 ltvoff=1.53357e-011               wtvoff=3.2331e-011 ptvoff=-2.15275e-018              kt1=-0.19390503                lkt1=3.1019883e-009 wkt1=-1.7199834e-009            pkt1=-2.6443803e-016            kt2=-0.081119383 wkt2=1.0732396e-009             ute=-1.2710103                 wute=5.3551437e-008 ua1=1.0428223e-009             lua1=-4.6414276e-017            wua1=-3.2428753e-017 pua1=3.4874435e-024             ub1=-8.7951553e-019            lub1=5.5793251e-026 wub1=1.7650088e-025             pub1=-1.0350741e-032            uc1=3.9283209e-010 luc1=-2.5732226e-018            wuc1=2.6139721e-018             puc1=-3.5887683e-025 at=60250.577                  jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-9.3988259e-011 pu0=2.9202309e-017             lvsat=0.00089799428              pvsat=8.3369419e-011 lpclm=3.0997244e-008             ppclm=-4.5347274e-015            wpdiblc2=-5.1734326e-010 ppdiblc2=3.628984e-017              laigbacc=1.472381e-010              paigbacc=-2.1520162e-017 lbigsd=2.4760012e-011             pbigsd=-5.1291714e-018            lkt2=9.9184296e-010 pkt2=-4.1412548e-017            lute=1.8391502e-008             pute=-4.0079207e-015 lat=-0.00081187248             leta0=1.6822863e-011             peta0=-4.6431102e-018 letab=2.2752285e-010             petab=-1.5058426e-017            wat=-0.0047078383 pat=3.7770836e-010             u0_ss=0.000680247                u0_ff=-0.000680247 wu0_ss=-1.87748e-10               wu0_ff=1.87748e-10                vsat_ss=-18882.7 vsat_ff=7250.05                    vsat_sf=7250.05                    vsat_fs=-4833.34 wvsat_ss=0.00215263                 wvsat_ff=1.1e-09                    wvsat_sf=1.1e-09 wvsat_fs=2.6e-10                    a0_ss=-0.850002                  a0_sf=-1.44815 a0_fs=0.850002                   la0_ss=7.39501e-08                la0_sf=1.25989e-07 la0_fs=-7.39501e-08               wa0_ss=1.1e-13                    wa0_sf=1.65089e-07 wa0_fs=-1.1e-13                   pa0_ss=3.3e-20                    pa0_sf=-1.43627e-14 pa0_fs=-3.3e-20                   pdiblc2_ss=-0.00405093                pdiblc2_fs=0.00405093 lpdiblc2_ss=1.30097e-10                lpdiblc2_fs=-1.30097e-10               lu0_ss=-3.46926e-11 lu0_ff=3.46926e-11                pu0_ss=9.57516e-18                pu0_ff=-9.57516e-18 lvsat_ss=0.00104991                 lvsat_ff=-0.00036975                lvsat_sf=-0.00036975 lvsat_fs=0.0002465                  pvsat_ss=-1.19689e-10               pvsat_ff=3.3e-17 pvsat_sf=3.3e-17                    pvsat_fs=-2.2e-17                   wpdiblc2_ss=7.04056e-10 wpdiblc2_fs=-7.04056e-10               ppdiblc2_ss=-3.59069e-17               ppdiblc2_fs=3.59069e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_mac.27 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.37170234 lvth0=-5.2961854e-010            wvth0=2.8674988e-009             pvth0=6.2441042e-017 k2=-0.031578608               lk2=-1.9343326e-009            wk2=1.1119656e-008 pk2=-3.1977196e-016            cit=-0.0070759444              lcit=4.7174297e-010 wcit=9.102442e-010              pcit=-3.7887441e-017            voff=-0.13033092 lvoff=-3.2692968e-009            wvoff=5.0328758e-009             pvoff=-1.6375953e-017 eta0=0.0076309373               weta0=-6.3413869e-010            etab=-0.025063581 wetab=1.2378745e-009             u0=0.013079189                wu0=8.4984393e-010 ua=-2.2704227e-009            lua=3.5723634e-017             wua=1.4290972e-016 pua=-5.0324348e-024            ub=2.1215294e-018             lub=-3.3265701e-026 wub=-6.191675e-026             pub=1.1713387e-033             uc=1.5908589e-010 luc=-6.9343574e-018            wuc=-2.1486781e-017            puc=7.986252e-025 vsat=67218.049                  wvsat=0.0011122508               a0=4.4102911 la0=-6.1512716e-007            wa0=-1.0263432e-006            pa0=8.6182592e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=0.2554496                  lketa=-2.0231939e-008 wketa=-9.8926683e-008            pketa=4.7814075e-015             pclm=0.62055728 wpclm=3.7578507e-008             pdiblc2=0.0012962963               ppdiblc2=0 lpdiblc2=0                          aigbacc=0.017867309                waigbacc=-5.1611318e-010 aigc=0.0060736294               laigc=-1.0418615e-011            waigc=-5.0338431e-012 paigc=2.0552048e-020             aigsd=0.0067518486               laigsd=-6.4154255e-011 waigsd=-1.6950532e-010            paigsd=7.2428184e-018             bigsd=0.0022414314 wbigsd=-2.3582397e-010            tvoff=0.0015315                  ltvoff=1.34511e-012 wtvoff=-6.43756e-011              ptvoff=2.77929e-018               kt1=-0.070490357 lkt1=-3.19216e-009              wkt1=-2.0344922e-008            pkt1=6.8543384e-016 kt2=-0.10096274                wkt2=1.9633924e-009             ute=-0.13185432 wute=-7.3888607e-008            ua1=1.5293824e-009             lua1=-7.1228839e-017 wua1=-1.1641171e-017            pua1=2.4272769e-024             ub1=-8.8240195e-019 lub1=5.5940458e-026             wub1=5.9483384e-026             pub1=-4.3828485e-033 uc1=8.7267807e-010             luc1=-2.7045368e-017            wuc1=-3.956462e-017 puc1=1.7922314e-024             at=-1103.0708                 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)' jtsswgd='1.5e-007*(1+0.55*iboffp_flag)'                                    lu0=-1.2151399e-011 pu0=-2.8701958e-017            lvsat=0.0014757176               pvsat=2.2546892e-010 lpclm=1.8900221e-008             ppclm=-3.1443964e-015            wpdiblc2=1.9422222e-010 laigbacc=-2.8916119e-010            paigbacc=2.0754975e-017             lbigsd=-8.6882517e-011 pbigsd=9.9046069e-018             lkt2=2.0038542e-009             pkt2=-8.6810341e-017 lute=-3.9705452e-008            pute=2.4915215e-015             lat=0.0023171635 leta0=1.5671109e-010             peta0=2.243574e-017              letab=9.6971944e-010 petab=-5.4827188e-017            wat=0.0019523611               pat=3.8038193e-011 u0_ss=-0.00252346                u0_ff=0.00093333                 wu0_ss=1.81274e-10 wu0_ff=7e-17                      vsat_ss=321.021                    vsat_ff=9333.3 vsat_sf=9333.3                     vsat_fs=-9333.3                    wvsat_ss=-0.00110059 wvsat_ff=7e-10                      wvsat_sf=7e-10                      wvsat_fs=-7e-10 a0_ss=-4.17037                   a0_ff=4.77037                    a0_sf=1.02222 a0_fs=4.17037                    la0_ss=2.43289e-07                la0_ff=-2.43289e-07 la0_sf=1.1e-13                    la0_fs=-2.43289e-07               wa0_ss=5.43818e-07 wa0_ff=-5.43822e-07               wa0_sf=-1.16534e-07               wa0_fs=-5.43818e-07 pa0_ss=-2.7735e-14                pa0_ff=2.77349e-14                pa0_sf=3.3e-20 pa0_fs=2.7735e-14                 pdiblc2_ss=-0.00150003                pdiblc2_fs=0.00150003 ppdiblc2_ss=-6.7e-23                   ppdiblc2_fs=6.7e-23                    lpdiblc2_ss=-2.2e-16 lpdiblc2_fs=2.2e-16                    at_ss=26271.6                    at_fs=16419.8 lu0_ss=1.28697e-10                lu0_ff=-4.76e-11                  pu0_ss=-9.24502e-18 pu0_ff=2.2e-24                    lvsat_ss=7.05185e-05                lvsat_ff=-0.000476 lvsat_sf=-0.000476                  lvsat_fs=0.000476                   pvsat_ss=4.62249e-11 pvsat_ff=2.2e-17                    pvsat_sf=2.2e-17                    pvsat_fs=-2.2e-17 wpdiblc2_ss=-8.9e-15                   wpdiblc2_fs=8.9e-15                    lat_ss=-0.00133985 lat_fs=-0.000837407               wat_ss=-0.00725096                wat_fs=-0.00453185 pat_ss=3.69799e-10                pat_fs=2.31124e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_mac.28 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.47365401 lvth0=3.7523517e-009             wvth0=9.0394144e-009             pvth0=-1.9677941e-016 k2=0.096477536                lk2=-7.3126906e-009            wk2=-1.1578264e-008 pk2=6.3354068e-016             cit=-0.011023377               lcit=6.3753513e-010 wcit=4.9875706e-010             pcit=-2.0604981e-017            voff=-0.21536309 lvoff=3.0205419e-010             wvoff=1.1790972e-008             pvoff=-3.0021599e-016 eta0=-0.0046404695              weta0=2.1514812e-009             etab=-0.018222363 wetab=1.9638846e-009             u0=0.014710738                wu0=1.0271143e-009 ua=-1.4826974e-009            lua=2.6391699e-018             wua=1.7998593e-017 pua=2.1383266e-025             ub=1.4789104e-018             lub=-6.2757053e-027 wub=9.9851737e-026             pub=-5.6229378e-033            uc=6.5843078e-011 luc=-3.0181593e-018            wuc=-1.8899121e-017            puc=6.8994351e-025 vsat=72071.205                  wvsat=0.011594661                a0=-1.1345781 la0=-3.8224265e-007            wa0=2.0359409e-006             pa0=-4.2433339e-014 ags=1                          lags=0                          wags=0 pags=0                          keta=-0.79692805                lketa=2.3967922e-008 wketa=6.7257402e-008             pketa=-2.1983241e-015            pclm=1.7478104 wpclm=-1.9703531e-007            pdiblc2=-0.0023703704              lpdiblc2=1.54e-010 aigbacc=0.015654395                waigbacc=-7.4264104e-010            aigc=0.0057959452 laigc=1.2441209e-012             waigc=-5.4431471e-012            paigc=3.7742812e-020 aigsd=0.0051882311               laigsd=1.51768e-012               waigsd=1.2944791e-011 paigsd=-4.2008638e-019            bigsd=0.0001728                  tvoff=0.00173375 ltvoff=-7.14943e-012              wtvoff=6.38928e-011               ptvoff=-2.60798e-018 kt1=-0.0019110449              lkt1=-6.0724911e-009            wkt1=-4.540691e-009 pkt1=2.1656137e-017             kt2=-0.086477086               wkt2=2.3398598e-009 ute=-0.74684197                wute=-7.1040015e-008            ua1=-8.28035e-010 lua1=2.7782691e-017             wua1=2.219837e-016              pua1=-7.3849678e-024 ub1=1.7867697e-018             lub1=-5.6164752e-026            wub1=-2.4920862e-025 pub1=8.5822157e-033             uc1=3.6282938e-010             luc1=-5.631723e-018 wuc1=3.798145e-017              puc1=-1.4647036e-024            at=18342.177 jtsswgs='1.5e-007*(1+0.55*iboffp_flag)'                                    jtsswgd='1.5e-007*(1+0.55*iboffp_flag)' lu0=-8.0676453e-011            pu0=-3.6147311e-017            lvsat=0.0012718851 pvsat=-2.1479231e-010            lpclm=-2.8444409e-008            ppclm=6.7093838e-015 wpdiblc2=1.9422222e-010             ppdiblc2=-9.9322927e-032            laigbacc=-1.9621881e-010 paigbacc=3.0269145e-017             lkt2=1.3954567e-009             pkt2=-1.0262197e-016 lute=-1.387597e-008             pute=2.3718806e-015             lat=0.0015004631 leta0=6.7211017e-010             peta0=-9.4560297e-017            letab=6.8238828e-010 petab=-8.531961e-017             wat=0.0015543808               pat=5.4753366e-011 cit_mc=0.0030963                  cit_mcl=-0.00495679                lcit_mc=-1.30044e-10 lcit_mcl=2.08185e-10                wcit_mc=-8.54578e-10               wcit_mcl=3.56074e-10 pcit_mc=3.58923e-17                pcit_mcl=-1.49551e-17               voff_ff=-0.0124938 voff_mc=-0.020642                  lvoff_ff=5.24741e-10                lvoff_mc=8.66963e-10 wvoff_ff=1.4243e-09                 wvoff_mc=5.69719e-09                pvoff_ff=-5.98204e-17 pvoff_mc=-2.39282e-16               eta0_mc=-0.00312346                weta0_mc=3.56074e-10 u0_ss=0.00252346                 u0_ff=-0.000308643               u0_sf=0.000733331 u0_fs=-0.000733331               wu0_ss=-1.81274e-10               wu0_ff=-7.12151e-11 wu0_sf=-3.7e-16                   wu0_fs=3.7e-16                    vsat_ss=-3160.46 vsat_ff=3160.46                    vsat_sf=-5666.7                    vsat_fs=5666.7 vsat_mc=4916.05                    wvsat_ss=0.0014243                  wvsat_ff=-0.0014243 wvsat_sf=-7e-10                     wvsat_fs=7e-10                      wvsat_mc=-0.00014243 a0_ss=7.57037                    a0_ff=-4.77037                   a0_sf=4.77037 a0_fs=-7.57037                   la0_ss=-2.49822e-07               la0_ff=1.57422e-07 la0_sf=-1.57422e-07               la0_fs=2.49822e-07                wa0_ss=-5.43818e-07 wa0_ff=5.43822e-07                wa0_sf=-5.43822e-07               wa0_fs=5.43818e-07 pa0_ss=1.79462e-14                pa0_ff=-1.79461e-14               pa0_sf=1.79461e-14 pa0_fs=-1.79462e-14               pdiblc2_ss=-0.00699997                pdiblc2_fs=0.00699997 lpdiblc2_ss=2.31e-10                   lpdiblc2_fs=-2.31e-10                  at_ss=4691.4 at_ff=-20642                     at_sf=-15481.5                   at_fs=4222.25 at_mc=-11000                     lu0_ss=-8.32739e-11               lu0_ff=4.56303e-12 lu0_sf=-3.08e-11                  lu0_fs=3.08e-11                   pu0_ss=5.98206e-18 pu0_ff=2.99102e-18                pu0_sf=-4.4e-24                   pu0_fs=4.4e-24 lvsat_ss=0.000216741                lvsat_ff=-0.000216741               lvsat_sf=0.000154 lvsat_fs=-0.000154                  lvsat_mc=-0.000206474               pvsat_ss=-5.98204e-11 pvsat_ff=5.98204e-11                pvsat_sf=-5.6e-17                   pvsat_fs=5.6e-17 pvsat_mc=5.98207e-12                wpdiblc2_ss=4.4e-15                    wpdiblc2_fs=-4.4e-15 ppdiblc2_ss=3.3e-23                    ppdiblc2_fs=-3.3e-23                   lat_ss=-0.000433477 lat_ff=0.000866963                lat_sf=0.000650222                lat_fs=-0.000325111 lat_mc=0.000462                   leta0_mc=1.31185e-10                peta0_mc=-1.49551e-17 wat_ss=-0.00129482                wat_ff=0.00569719                 wat_sf=0.00427289 wat_fs=-0.00116534                wat_mc=4.4e-09                    pat_ss=1.19641e-10 pat_ff=-2.39282e-10               pat_sf=-1.79461e-10               pat_fs=8.97309e-11 pat_mc=3.3e-17 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_12_mac.global nmos ( modelid=7                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_12'              permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=2.42e-009                  toxm=2.42e-009                  dtox=2.4017e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=-1.2e-008 xw=6e-009                     dlc=7.5e-009                   dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.42161 k3=-6.68                      k3b=0.645                      w0=0 dvt0=0.13719                    dvt1=0.37921                    dvt2=-0.1 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.60407                    minv=-0.5                       voffl=0 dvtp0=4.2e-007                   dvtp1=5                          lpe0=1e-009 lpeb=0                          xj=6.7e-008                   ngate=3e+021 ndep=1e+017                     nsd=1e+020                     phin=0.13 cdsc=0                          ud=0                          cdscb=0 cdscd=0                          nfactor=0.7                        a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=1                          drout=0.56                       pvag=2 delta=0.01                       pscbe1=1e+009                     pscbe2=1e-020 fprout=0                          pdits=0.0025                     pditsd=0.99219 pditsl=0                          rsh=18                         rdsw=111.62 prwg=0                          prwb=0                          wr=1 alpha0=1e-008                     alpha1=0.3                        beta0=11.7 bgidl=2.5e+008                   cgidl=12.928                     egidl=0.17539 bigbacc=0.0054245                  cigbacc=0.2809                     nigbacc=3.5692851 aigbinv=0.013093326                bigbinv=0.0028088446               cigbinv=0.006 eigbinv=1.1                        nigbinv=2.6384376                  bigc=0.0011209 cigc=1e-005                     bigsd=0.00059897493              cigsd=2e-020 nigc=2.3705874                  poxedge=1                          pigcd=2.2301237 ntox=1                          vfbsdoff=0.01                       cgso=1e-010 cgdo=1e-010                     cgbo=0                          cgdl=5e-012 cgsl=5e-012                     clc=0                          cle=0.6 cf='6.7e-011+9.3e-011*ccoflag_12'                                     ckappas=0.6 ckappad=0.6                        acde=0.3                        moin=5 noff=2.7                        voffcv=-0.16                      tvfbsdoff=0.01015 kt1l=0                          prt=0                          fnoimod=1.000000e+00 tnoimod=0                          em=1.000000e+06               ef=8.500000e-01 noia=0                          noib=0                          noic=0 jss=2.24e-07                   jsd=2.24e-07                   jsws=7.31e-14 jswd=7.31e-14                   jswgs=7.31e-14                   jswgd=7.31e-14 njs=1.02                       njd=1.02                       ijthsfwd=0.01 ijthdfwd=0.01                       ijthsrev=0.01                       ijthdrev=0.01 bvs=8.22                       bvd=8.22                       xjbvs=1 xjbvd=1                          njtsswg=10                         xtsswgs=0.31 xtsswgd=0.31                       tnjtsswg=0.5                        vtsswgs=8 vtsswgd=8                          pbs=0.672                      pbd=0.672 cjs=0.00144                    cjd=0.00144                    mjs=0.327 mjd=0.327                      pbsws=0.438                      pbswd=0.438 cjsws=1.13e-010                  cjswd=1.13e-010                  mjsws=0.008 mjswd=0.008                      pbswgs=0.9                        pbswgd=0.9 cjswgs=2.7e-010                   cjswgd=2.7e-010                   mjswgs=0.779 mjswgd=0.779                      tpb=0.0013                     tcj=0.0008 tpbsw=0.00218                    tcjsw=0.00016                    tpbswg=0.0012 tcjswg=0.00107                    xtis=3                          xtid=3 dmcg=4.2e-008                   dmci=4.2e-008                   dmdg=0 dmcgt=0                          dwj=0                          xgw=0 xgl=2.64e-009                  rshg=16.42                      gbmin=1e-012 rbpb=50                         rbpd=50                         rbps=50 rbdb=50                         rbsb=50                         ngcon=1 xrcrg1=12                         xrcrg2=1                          k2we=0 ku0we=-0.0018                    kvth0we=0.0010                     lk2we=0e-11 lku0we=9e-12                      lkvth0we=-3e-011                    pk2we=0e-18 pku0we=0e-17                      pkvth0we=2.5e-018                   scref=1e-6 web=1251.3                     wec=-6544.5                    wk2we=0e-11 wku0we=3e-11                      wkvth0we=-7e-011                    wpemod=1 lintnoi=-5e-08 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.11 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.6 iboffn_flag='iboffn_flag_12' iboffp_flag='iboffp_flag_12' sigma_factor='sigma_factor_12' ccoflag='ccoflag_12' rcoflag='rcoflag_12' rgflag='rgflag_12' mismatchflag='mismatchflag_mos_12' globalflag='globalflag_mos_12' totalflag='totalflag_mos_12' global_factor='global_factor_12' local_factor='local_factor_12' sigma_factor_flicker='sigma_factor_flicker_12' noiseflag='noiseflagn_12' noiseflag_mc='noiseflagn_12_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w1='2.3875*0.35355' w2='0.70711*-0.35355' w3='0.54772*-0.0052117' w4='0.54772*-0.40307' w5='0.54772*-0.64548' w6='0.54772*-0.049915' w7='0.54772*-0.11513' w8='0.54772*-0.39385' w9='0' w10='0' tox_c='toxn_12'                  dxl_c='dxln_12'                  dxw_c='dxwn_12' cj_c='cjn_12'                   cjsw_c='cjswn_12'                 cjswg_c='cjswgn_12' cgo_c='cgon_12'                  cgl_c='cgln_12'                  ddlc_c='ddlcn_12' ntox_c='ntoxn_12'                 cf_c='cfn_12'                   dvth_c='dvthn_12' dlvth_c='dlvthn_12'                dwvth_c='dwvthn_12'                dpvth_c='dpvthn_12' du0_c='du0n_12'                  dlu0_c='dlu0n_12'                 dwu0_c='dwu0n_12' dpu0_c='dpu0n_12'                 dvsat_c='dvsatn_12'                dlvsat_c='dlvsatn_12' dwvsat_c='dwvsatn_12'               dpvsat_c='dpvsatn_12'               dk2_c='dk2n_12' dlk2_c='dlk2n_12'                 dwk2_c='dwk2n_12'                 dpk2_c='dpk2n_12' dags_c='dagsn_12'                 dlags_c='dlagsn_12'                dwags_c='dwagsn_12' dpags_c='dpagsn_12'                dcit_c='dcitn_12'                 dlcit_c='dlcitn_12' dwcit_c='dwcitn_12'                dpcit_c='dpcitn_12'                dpclm_c='dpclmn_12' dlpclm_c='dlpclmn_12'               dwpclm_c='dwpclmn_12'               dppclm_c='dppclmn_12' dua1_c='dua1n_12'                 dlua1_c='dlua1n_12'                dwua1_c='dwua1n_12' dpua1_c='dpua1n_12'                duc_c='ducn_12'                  dluc_c='dlucn_12' dwuc_c='dwucn_12'                 dpuc_c='dpucn_12'                 dketa_c='dketan_12' dlketa_c='dlketan_12'               dwketa_c='dwketan_12'               dpketa_c='dpketan_12' jtsswg_c='jtsswgn_12'               ss_flag_c='ss_flagn_12'              ff_flag_c='ff_flagn_12' sf_flag_c='sf_flagn_12'              fs_flag_c='fs_flagn_12'              monte_flag_c='monte_flagn_12' c1f_c='c1fn_12'                  c2f_c='c2fn_12'                  c3f_c='c3fn_12' global_mc='global_mc_flag_12' tox_g='toxn_12_ms_global'        dxl_g='dxln_12_ms_global'        dxw_g='dxwn_12_ms_global' cj_g='cjn_12_ms_global'         cjsw_g='cjswn_12_ms_global'       cjswg_g='cjswgn_12_ms_global' cgo_g='cgon_12_ms_global'        cgl_g='cgln_12_ms_global'        ntox_g='ntoxn_12_ms_global' cf_g='cfn_12_ms_global'         dvth_g='dvthn_12_ms_global'       dlvth_g='dlvthn_12_ms_global' dwvth_g='dwvthn_12_ms_global'      dpvth_g='dpvthn_12_ms_global'      du0_g='du0n_12_ms_global' dlu0_g='dlu0n_12_ms_global'       dwu0_g='dwu0n_12_ms_global'       dpu0_g='dpu0n_12_ms_global' dvsat_g='dvsatn_12_ms_global'      dlvsat_g='dlvsatn_12_ms_global' dwvsat_g='dwvsatn_12_ms_global'     dpvsat_g='dpvsatn_12_ms_global'     dk2_g='dk2n_12_ms_global' dlk2_g='dlk2n_12_ms_global'       dwk2_g='dwk2n_12_ms_global'       dpk2_g='dpk2n_12_ms_global' dags_g='dagsn_12_ms_global'       dwags_g='dwagsn_12_ms_global'      dcit_g='dcitn_12_ms_global' dlcit_g='dlcitn_12_ms_global'      dwcit_g='dwcitn_12_ms_global'      dpcit_g='dpcitn_12_ms_global' dpclm_g='dpclmn_12_ms_global'      dlpclm_g='dlpclmn_12_ms_global' dwpclm_g='dwpclmn_12_ms_global'     dpua1_g='dpua1n_12_ms_global'      dluc_g='dlucn_12_ms_global' dlketa_g='dlketan_12_ms_global'     dwketa_g='dwketan_12_ms_global' ss_flag_g='ss_flagn_12_ms_global'    ff_flag_g='ff_flagn_12_ms_global' monte_flag_g='monte_flagn_12_ms_global'                                        sf_flag_g='sf_flagn_12_ms_global' fs_flag_g='fs_flagn_12_ms_global' weight1=-3.3988235 weight2=2.0543791 weight3=1.2109804 weight4=-0.65359477 weight5=-0.4543268 tox_1=4.3370683e-012 tox_2=-9.3347319e-012 tox_3=-3.153177e-012 tox_4=3.7476726e-011 tox_5=7.3686462e-013 dxl_1=2.1275845e-010 dxl_2=-4.5792666e-010 dxl_3=-1.5467887e-010 dxl_4=-1.8384866e-009 dxl_5=3.6147736e-011 dxw_1=-6.4604528e-010 dxw_2=-8.7924358e-010 dxw_3=2.9521784e-010 dxw_4=-2.4998818e-025 dxw_5=-5.892057e-009 cj_1=9.4508e-006 cj_2=-1.865e-006 cj_3=-5.1171e-006 cj_4=-6.1145e-021 cj_5=-1.0203e-006 cjsw_1=7.4162e-013 cjsw_2=-1.4635e-013 cjsw_3=-4.0155e-013 cjsw_4=-8.8584e-028 cjsw_5=-8.0062e-014 cjswg_1=1.772e-012 cjswg_2=-3.4968e-013 cjswg_3=-9.5946e-013 cjswg_4=-2.1166e-027 cjswg_5=-1.913e-013 cgo_1=-6.563e-013 cgo_2=1.2951e-013 cgo_3=3.5536e-013 cgo_4=7.8393e-028 cgo_5=7.0851e-014 cgl_1=-3.2815e-014 cgl_2=6.4755e-015 cgl_3=1.7768e-014 cgl_4=8.2778e-029 cgl_5=3.5426e-015 ntox_1=-0.14705 ntox_2=0.026969 ntox_3=0.18642 ntox_4=3.0066e-016 ntox_5=0.021676 cf_1=-4.3972e-013 cf_2=8.6772e-014 cf_3=2.3809e-013 cf_4=5.3077e-028 cf_5=4.747e-014 dvth_1=0.0021309 dvth_2=0.0040543 dvth_3=-0.00048665 dvth_4=2.4146e-018 dvth_5=-0.00085354 dlvth_1=1.0938e-010 dlvth_2=3.6124e-011 dlvth_3=-5.9806e-011 dlvth_4=1.4564e-025 dlvth_5=-2.0322e-011 dwvth_1=3.0174e-010 dwvth_2=6.7977e-011 dwvth_3=-1.2704e-010 dwvth_4=7.1369e-025 dwvth_5=-4.9451e-011 dpvth_1=2.4461e-017 dpvth_2=8.7501e-018 dpvth_3=-1.332e-017 dpvth_4=1.7894e-032 dpvth_5=-4.4473e-018 du0_1=4.9704e-005 du0_2=0.00028611 du0_3=8.7773e-006 du0_4=1.8414e-020 du0_5=-4.876e-005 dlu0_1=-6.5208e-012 dlu0_2=1.6953e-011 dlu0_3=5.7318e-012 dlu0_4=1.4918e-026 dlu0_5=-1.5045e-012 dwu0_1=1.1013e-011 dwu0_2=1.8005e-011 dwu0_3=-1.2862e-012 dwu0_4=-8.9741e-027 dwu0_5=-3.9519e-012 dpu0_1=-1.0722e-018 dpu0_2=2.272e-018 dpu0_3=1.0589e-018 dpu0_4=1.4779e-033 dpu0_5=-2.4256e-019 dvsat_1=103.72 dvsat_2=1340.2 dvsat_3=110.4 dvsat_4=-1.4859e-013 dvsat_5=-209.11 dlvsat_1=2.3813e-005 dlvsat_2=4.3272e-005 dlvsat_3=-7.1286e-006 dlvsat_4=-2.2296e-021 dlvsat_5=-9.3263e-006 dwvsat_1=1.1926e-005 dwvsat_2=0.00015763 dwvsat_3=8.7283e-006 dwvsat_4=-6.1118e-020 dwvsat_5=-2.4025e-005 dpvsat_1=4.2356e-012 dpvsat_2=1.0453e-011 dpvsat_3=-5.9474e-012 dpvsat_4=-1.845e-026 dpvsat_5=-2.3051e-012 dk2_1=0.0032033 dk2_2=-0.00063675 dk2_3=-0.0014925 dk2_4=1.7091e-018 dk2_5=-0.00033267 dlk2_1=4.6723e-011 dlk2_2=1.8218e-010 dlk2_3=2.3162e-011 dlk2_4=-8.4614e-027 dlk2_5=-3.0686e-011 dwk2_1=5.8553e-012 dwk2_2=-1.3642e-012 dwk2_3=7.7152e-012 dwk2_4=3.0896e-027 dwk2_5=-4.0857e-014 dpk2_1=-1.6392e-018 dpk2_2=3.9307e-019 dpk2_3=-2.741e-018 dpk2_4=-5.206e-033 dpk2_5=-2.012e-020 dags_1=0.017847 dags_2=0.0207 dags_3=0.0099509 dags_4=1.3481e-018 dags_5=-0.0044963 dwags_1=-9.7014e-010 dwags_2=6.3029e-010 dwags_3=-1.6335e-010 dwags_4=-1.307e-024 dwags_5=5.5423e-011 dcit_1=2.5697e-006 dcit_2=-5.7337e-007 dcit_3=2.0649e-006 dcit_4=1.9353e-021 dcit_5=-8.9683e-008 dlcit_1=-2.2774e-012 dlcit_2=5.0797e-013 dlcit_3=-1.8203e-012 dlcit_4=-2.3229e-028 dlcit_5=8.0013e-014 dwcit_1=-2.3201e-013 dwcit_2=4.9456e-014 dwcit_3=-6.5829e-014 dwcit_4=-1.8151e-028 dwcit_5=1.4648e-014 dpcit_1=2.0574e-019 dpcit_2=-4.3833e-020 dpcit_3=5.7145e-020 dpcit_4=4.641e-035 dpcit_5=-1.3057e-020 dpclm_1=-0.011251 dpclm_2=0.0022202 dpclm_3=0.0060918 dpclm_4=1.5339e-017 dpclm_5=0.0012146 dlpclm_1=-1.4064e-009 dlpclm_2=2.7752e-010 dlpclm_3=7.6148e-010 dlpclm_4=-4.5358e-025 dlpclm_5=1.5182e-010 dwpclm_1=-1.1332e-009 dwpclm_2=2.1201e-010 dwpclm_3=1.2183e-009 dwpclm_4=-8.462e-025 dwpclm_5=1.5518e-010 dpua1_1=-1.0928e-026 dpua1_2=2.6204e-027 dpua1_3=-1.8273e-026 dpua1_4=2.1063e-042 dpua1_5=-1.3413e-028 dluc_1=1.6392e-020 dluc_2=-3.9307e-021 dluc_3=2.741e-020 dluc_4=-2.049e-035 dluc_5=2.012e-022 dlketa_1=-4.3713e-010 dlketa_2=1.0482e-010 dlketa_3=-7.3092e-010 dlketa_4=-7.9139e-025 dlketa_5=-5.3653e-012 dwketa_1=-1.6392e-010 dwketa_2=3.9307e-011 dwketa_3=-2.741e-010 dwketa_4=-1.2123e-026 dwketa_5=-2.012e-012 ss_flag_1=0.039117 ss_flag_2=-0.0053993 ss_flag_3=-0.14213 ss_flag_4=1.7869e-016 ss_flag_5=-0.010792 ff_flag_1=-0.054641 ff_flag_2=0.013102 ff_flag_3=-0.091365 ff_flag_4=3.509e-017 ff_flag_5=-0.00067066 monte_flag_1=0.0818308 monte_flag_2=-0.176127 monte_flag_3=-0.0594923 monte_flag_4=-0.707115 monte_flag_5=0.0139031 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.98 b_4=-0.009                     c_4=-0.012                     d_4=0.0005 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.0031                     mis_a_2=0.15                       mis_a_3=-0.15 mis_b_1=0.0030                     mis_b_2=-0.05                      mis_b_3=0.08 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.00083                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.0035                     mis_e_2=0.05                       mis_e_3=0.03 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-1.2e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18                         bidirectionflag=1 designflag=1 cf0=6.7e-011                   cco=9.3e-011 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=1.0                        l_rjtsswg=0                          ll_rjtsswg=2 w_rjtsswg=0.0e-03                    ww_rjtsswg=2                          p_rjtsswg=0 noimod=1                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6                sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=0                   lreflod=1e-6                llodref=3 lod_clamp=-1e-90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=0 kvth00=0                   lkvth00=0                   wkvth00=0 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=0                   lku000=0                   wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0                   lkvth000=0                   wkvth000=0         		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=-6e-2                   wku01=0 pku01=0                   llodku01=-1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=3e-2                   wkvth01=0 pkvth01=0                   llodvth1=-1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.00               lku02=0e-7              wku02=0e-8 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0.9 kvth02=0e-3                lkvth02=0e-9               wkvth02=0e-9 pkvth02=0e-15               llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=-0e-2 lodeta02=1 wlod02=0 ku002=-0.050                   lku002=17e-10                  wku002=18e-10	           pku002=-11e-17 llodku002=1                   wlodku002=1 kvth002=-9e-3                   lkvth002=6.7e-10                  wkvth002=13e-10                 pkvth002=-5.5e-17 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=-0.0              lku03=-0e-9               wku03=-0e-8 pku03=0e-15                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0.3 kvth03=0e-3                lkvth03=-0e-9               wkvth03=-0e-8 pkvth03=-0e-16               llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=-0.028                   lku003=-1e-10                  wku003=-5.5e-9	           pku003=-7e-17 llodku003=1                   wlodku003=1 kvth003=-2e-3                   lkvth003=5e-10                  wkvth003=8e-10                 pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=0.991e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=10.01e-6                w_b1=10e-6 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=-0.5e-8              wdpcku0=1 lku0dpc=-0.1e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=-6                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='0.10'              wkvth0dpl=0                   wdplkvth0=1 lkvth0dpl='3.0e-8*1*1.5'              ldplkvth0=1.0                 pkvth0dpl=0 ku0dpl=' 0.7*1+0.1'                wku0dpl='1e-8*0'                   wdplku0=1 lku0dpl='2.8e-5*1'              ldplku0=0.7                 pku0dpl=1e-14 keta0dpl='0.2'                wketa0dpl=0                   wdplketa0=1 kvsatdpl='0.5*0'                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx=0.0                wku0dpx=0e-9                wdpxku0=1 lku0dpx=0.0e-8              ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=0.02               wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-2             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='0.0'               wku0dps=0                   wdpsku0=1 lku0dps='0e-8'             ldpsku0=1.0                 pku0dps=0 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0.0                 wdps=0 kvth0dps_b1=-0.00            kvth0dps_b2=-0.000            dpsbinflg=1 ku0dps_b1=0.0                ku0dps_b2=0.04 keta0dps_b1=0                  keta0dps_b2=0.02 kvth0dpa='0.055'               wkvth0dpa=-0.0e-9            wdpakvth0=1 lkvth0dpa=0.001e-7            ldpakvth0=1.0                pkvth0dpa=-0.0e-17 ku0dpa='0.18'               wku0dpa=0e-9               wdpaku0=1 lku0dpa=1e-9               ldpaku0=1.0                 pku0dpa=5e-16 keta0dpa=0.035                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0.6                wdpa=0 kvth0dpa_b1=0             kvth0dpa_b2=0.04            dpabinflg=1 ku0dpa_b1=-0.00             ku0dpa_b2=0.035 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2=0.012               wkvth0dp2=0.2e-8             wdp2kvth0=1 lkvth0dp2='2.0e-9*1.5'              ldp2kvth0=1.0                   pkvth0dp2=0 ku0dp2='0.03'                wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2='2.5e-7'              ldp2ku0=0.7                 pku0dp2=0 keta0dp2='0.01*0'                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=1.5                wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.05            kvth0dp2l_b2=0.00           dp2lbinflg=1 ku0dp2l_b1='-0.03'            ku0dp2l_b2=0.0 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a='0.05'              wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a='1.0e-9*0'             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.1              wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=4.0e-8            ldp2aku0=1.0                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.05               wdp2a=0 kvth0dp2a_b1=0.00           kvth0dp2a_b2=0.05           dp2abinflg=1 ku0dp2a_b1=0.24                ku0dp2a_b2=0.05 keta0dp2a_b1=0.0                 keta0dp2a_b2=0.02 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5     enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx=0.03                wkvth0enx='3.0e-9'            wenxkvth0=1.0 lkvth0enx='-11.0e-9*0'        lenxkvth0=1.0                 pkvth0enx='6e-16' ku0enx=-1.0                wku0enx='-5.0e-8'    wenxku0=1.0 lku0enx=1.5e-8              lenxku0=1.2                 pku0enx='4.5e-17' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx='1.0*0'             wka0enx='1e-6*0'            wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx='1.2'               wenx=0                   ku0enx0='-0.20*0' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.05e-6 kvth0eny='0.010*5'           wkvth0eny='1.0e-9*2.0'        wenykvth0=1 lkvth0eny='1.0e-7*1.5'        lenykvth0=1.0                 pkvth0eny=0 ku0eny='-0.30-0.1'         wku0eny=-1.5e-8             wenyku0=1 ku0eny0='-0.01*2.0'         wku0eny0='-1.0e-7*1.0'       weny0ku0=1 lku0eny='3.0e-10+2.0e-10'   lenyku0=1.5                 pku0eny='0.9e-19*1' keta0eny=0e-4                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny='0.7'               weny=0 kvth0eny1='-6e-4*1'          wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1='3.0e-18*1' ku0eny1='0.003*0'          wku0eny1='-1.0e-10*0'       weny1ku0=1 lku0eny1='0.6e-8*0'         leny1ku0=1.0                pku0eny1='-5.5e-17*0' keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1='1.0e-8*0'         weny1ka0=1 lka0eny1='4.0e-9*0'         leny1ka0=1.0                pka0eny1='3.0e-15*0' kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5              ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=-0.036              wkvth0rx=-4.0e-9             wrxkvth0=1.0 lkvth0rx=2.3e-08             lrxkvth0=1.0                 pkvth0rx=-2.5e-16 ku0rx=0.5                 wku0rx=5.2e-8              wrxku0=1.0 lku0rx=5e-10             lrxku0=1.2                 pku0rx=0.0e-17 keta0rx=0.0                 wketa0rx=0                   wrxketa0=1 kvsatrx=0.5                 wrx=0                   ku0rx0=-0.1 ry_mode=1 ringymax=0.9027e-5           ringymin=0.117e-6 ryref=1.8027e-5 kvth0ry=-0.04               wkvth0ry=-3.0e-9             wrykvth0=1.0 lkvth0ry=0.0e-8               lrykvth0=1.0                 pkvth0ry=-2.5e-16 ku0ry=0.170                wku0ry=5.0e-8              wryku0=1.0 lku0ry=0.8e-9               lryku0=1.1                 pku0ry=-0.0e-17 keta0ry=0.00                 wketa0ry=0                   wryketa0=1 kvsatry=0.2                  wry=0 kvth0ry0=-0.0                 ku0ry0=0.0 sfxref=9.0e-8            sfxmax=3.906e-6           minwodx=0.0e-6 sfxmin=9.0e-8 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a='-0.000'            lkvth0odx1a='1.0e-13*0'           lodx1akvth0='2.0' wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.90 kvth0odx1b=-0.0009           lkvth0odx1b='0+3e-12-1e-12'            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b='-0.0028-0.0005'           lku0odx1b=1e-10           lodx1bku0=1.0 wku0odx1b=-0.8e-10          wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6 sfymax=10e-6             minwody=0.9e-6            wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-0.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.2 lrefody=5e-8              lodyref=1 kvth0odyb=0.018             lkvth0odyb=-8.0e-10          lodybkvth0=1.0 wkvth0odyb=-10.5e-8          wodybkvth0=1.0               pkvth0odyb=-0.5e-15 ku0odyb=0.01              lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-0.5e-7           wodybku0=1.0               pku0odyb=0.2e-15 web_mac=2153.1  wec_mac=-9093.6 kvsatwe=0.0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_12_mac.1 nmos ( level=54                         lmin=9e-007                     lmax=9.019e-06 wmin=9e-007                     wmax=9.007e-06                  vth0=0.47770481 lvth0=1.3593445e-008             wvth0=-4.4942852e-009            pvth0=9.5709661e-016 k2=-0.012512956               lk2=-2.4224835e-009            wk2=-1.5154349e-008 pk2=3.2176839e-016             cit=0.0024988694               lcit=-4.3033167e-010 wcit=-7.9574053e-011            pcit=4.7982407e-017             voff=-0.1867703 lvoff=-1.1897818e-008            wvoff=-1.225929e-008             pvoff=1.0430929e-015 eta0=0.0094474074               weta0=-4.0293511e-009            etab=-0.050049327 wetab=4.4423596e-010             u0=0.019440236                lu0=2.1323393e-009 wu0=2.7607987e-009             pu0=5.6416838e-016             ua=-1.3720449e-009 lua=1.2741052e-017             wua=1.2162378e-016             pua=2.7778165e-023 ub=1.679841e-018              lub=1.1232431e-025             wub=7.4216595e-026 pub=-4.6863043e-032            uc=9.871264e-011              luc=1.9416514e-017 wuc=-5.428261e-018             puc=-1.0342625e-023            vsat=100000 a0=1.241187                   la0=7.0366792e-007             wa0=9.2887001e-008 pa0=2.644477e-014              ags=0.45083774                 lags=6.2323126e-007 wags=6.7013754e-008             pags=-1.3879161e-014            keta=-0.012870078 lketa=-4.3467431e-008            wketa=1.6003697e-008             pketa=3.4295672e-016 pclm=1.1419915                  lpclm=2.1714219e-008             wpclm=2.2758372e-008 ppclm=2.4814535e-013             pdiblc2=0.0011708574               lpdiblc2=2.3615201e-009 wpdiblc2=-2.7329357e-010            ppdiblc2=1.4111136e-015             agidl=2.0002496e-010 lagidl=-2.1526588e-017            wagidl=-4.3823313e-017            pagidl=1.5116522e-023 aigbacc=0.013531                   aigc=0.011455023                laigc=-3.9097721e-011 waigc=-2.3988795e-011            paigc=-3.3404334e-018            aigsd=0.010832691 laigsd=-4.3085085e-012            waigsd=5.9855909e-012             paigsd=4.6743834e-017 tvoff=0.00205632                 ltvoff=-2.80529e-011              wtvoff=-2.37966e-010 ptvoff=-4.35451e-017              kt1=-0.15041256                lkt1=-6.0675673e-009 wkt1=5.1763833e-009             pkt1=6.5375977e-016             kt2=-0.068219259 lkt2=1.9707022e-009             ute=-0.69752755                lute=-1.3155948e-008 wute=-8.1480464e-008            pute=8.2453737e-014             ua1=1.6294632e-009 lua1=-1.8024572e-016            wua1=-9.5584212e-017            pua1=1.4130996e-022 ub1=-9.4068388e-019            lub1=2.0665324e-025             wub1=1.4079127e-025 pub1=-6.243337e-032             uc1=2.5354731e-010             luc1=3.7650631e-017 wuc1=5.4643971e-017             puc1=1.5881302e-023             at=121006.13 lat=-0.0090431364              wat=0.00063308461              pat=-5.6901644e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' lvsat=0                          wvsat=0                          pvsat=0 ags_ff=0.112177                   ags_ss=-0.112177                  ags_fs=0.0899896 ags_sf=-0.0788959                 lags_ff=-9.96137e-08               lags_ss=9.96137e-08 lags_fs=-7.99108e-08               lags_sf=7.00595e-08                wags_ff=-1.11745e-08 wags_ss=1.11745e-08                wags_fs=-1.11742e-08               wags_sf=1.11741e-08 pags_ff=9.92269e-15                pags_ss=-9.92269e-15               pags_fs=9.9227e-15 pags_sf=-9.92266e-15 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_12_mac.2 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=9.007e-06                  vth0=0.48875521 lvth0=3.780688e-009              wvth0=-2.0212307e-009            pvth0=-1.2389758e-015 k2=-0.015187625               lk2=-4.7377755e-011            wk2=-1.4102816e-008 pk2=-6.1199289e-016            cit=0.001871605                lcit=1.266791e-010 wcit=-2.2044158e-010            pcit=1.7307277e-016             voff=-0.19131842 lvoff=-7.8590871e-009            wvoff=-1.3946656e-008            pvoff=2.5414734e-015 eta0=0.0094474074               weta0=-4.0293511e-009            etab=-0.050049327 wetab=4.4423596e-010             u0=0.020804506                lu0=9.2086745e-010 wu0=5.3180269e-009             pu0=-1.7066502e-015            ua=-1.4202214e-009 lua=5.5521798e-017             wua=2.9108738e-016             pua=-1.2270551e-022 ub=1.9446717e-018             lub=-1.2284538e-025            wub=1.6654941e-026 pub=4.2517047e-033             uc=1.3444957e-010             luc=-1.2317877e-017 wuc=2.8188979e-018             puc=-1.7666102e-023            vsat=100000 a0=2.2168401                  la0=-1.6271207e-007            wa0=1.2364369e-007 pa0=-8.6717083e-016            ags=0.9215647                  lags=2.0522571e-007 wags=1.3748303e-007             pags=-7.6455877e-014            keta=-0.042260195 lketa=-1.7369008e-008            wketa=1.5552113e-008             pketa=7.4396343e-016 pclm=1.0582242                  lpclm=9.6099579e-008             wpclm=4.0024888e-007 ppclm=-8.7066219e-014            pdiblc2=0.0043431329               lpdiblc2=-4.5546051e-010 wpdiblc2=1.5297986e-009             ppdiblc2=-1.9003217e-016            agidl=2.0166125e-010 lagidl=-2.2979613e-017            wagidl=-4.2121133e-017            pagidl=1.3604986e-023 aigbacc=0.013531                   aigc=0.01144156                 laigc=-2.7142719e-011 waigc=-2.7924578e-011            paigc=1.5454254e-019             aigsd=0.010901812 laigsd=-6.5688064e-011            waigsd=1.1012432e-010             paigsd=-4.5731357e-017 tvoff=0.00210505                 ltvoff=-7.13234e-011              wtvoff=-1.78508e-010 ptvoff=-9.63437e-017              kt1=-0.15829663                lkt1=9.3348849e-010 wkt1=2.04908e-008               pkt1=-1.2945443e-014            kt2=-0.079408928 lkt2=1.1907128e-008             ute=-0.7148261                 lute=2.2051684e-009 wute=2.6374118e-008             pute=-1.3321132e-014            ua1=1.8577961e-009 lua1=-3.8300532e-016            wua1=-2.2869608e-016            pua1=2.595133e-022 ub1=-1.1416261e-018            lub1=3.8508993e-025             wub1=5.5410293e-025 pub1=-4.2945412e-031            uc1=3.2268666e-010             luc1=-2.3745111e-017 wuc1=1.8234157e-016             puc1=-9.7514165e-023            at=173114.6 lat=-0.055315449               wat=-0.017369901               pat=1.0296486e-008 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-1.9609509e-009            pkt2=1.7413244e-015             lvsat=0 wvsat=0                          pvsat=0                          vsat_ff=5840 vsat_ss=-5948.77                   lvsat_ff=-0.00518592                lvsat_ss=0.00528251 wvsat_ff=1.6e-09                    wvsat_ss=0.000980389                pvsat_ff=6e-16 pvsat_ss=-8.70587e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_12_mac.3 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=9.007e-06                  vth0=0.50299904 lvth0=-2.4581081e-009            wvth0=-2.0323861e-010            pvth0=-2.0352563e-015 k2=-0.020631836               lk2=2.3371869e-009             wk2=-1.2542381e-008 pk2=-1.2954633e-015            cit=0.0021101629               lcit=2.2190745e-011 wcit=-4.3607509e-011            pcit=9.5619449e-017             voff=-0.19960549 lvoff=-4.2293521e-009            wvoff=-1.8136349e-008            pvoff=4.376559e-015 eta0=0.0094474074               weta0=-4.0293511e-009            etab=-0.050049327 wetab=4.4423596e-010             u0=0.022392389                lu0=2.2537489e-010 wu0=3.0812091e-009             pu0=-7.2692405e-016            ua=-1.290679e-009 lua=-1.2177874e-018            wua=4.8984204e-017             pua=-1.6664323e-023 ub=1.8293472e-018             lub=-7.2333239e-026            wub=8.5102635e-026 pub=-2.5728385e-032            uc=1.2753024e-010             luc=-9.287213e-018 wuc=-2.3074647e-017            puc=-6.3247295e-024            vsat=102729.69 a0=2.3695594                  la0=-2.2960313e-007            wa0=4.6874792e-007 pa0=-1.5202282e-013            ags=1.7828746                  lags=-1.7202802e-007 wags=-5.4361812e-007            pags=2.2186643e-013             keta=-0.038045373 lketa=-1.92151e-008              wketa=1.4725858e-008             pketa=1.1058632e-015 pclm=1.0886439                  lpclm=8.2775761e-008             wpclm=3.3319634e-007 ppclm=-5.7697208e-014            pdiblc2=0.0010595861               lpdiblc2=9.8273299e-010 wpdiblc2=-1.0667953e-010            ppdiblc2=5.2674524e-016             agidl=1.521082e-010 lagidl=-1.2753756e-018            wagidl=-9.2842719e-018            pagidl=-7.7755874e-025 aigbacc=0.013531                   aigc=0.011401792                laigc=-9.7244857e-012 waigc=-5.3328408e-011            paigc=1.128142e-017              aigsd=0.010750421 laigsd=6.2120975e-013             waigsd=-1.7149512e-011            paigsd=1.0014581e-017 tvoff=0.00207493                 ltvoff=-5.81302e-011              wtvoff=-4.42325e-010 ptvoff=1.92079e-017               kt1=-0.14221842                lkt1=-6.1087684e-009 wkt1=-1.3870336e-008            pkt1=2.1047353e-015             kt2=-0.050480114 lkt2=-7.6369231e-010            ute=-0.7401225                 lute=1.3284991e-008 wute=-7.560974e-009             pute=1.5424387e-015             ua1=8.9427012e-010 lua1=3.9019048e-017             wua1=7.1927351e-016             pua1=-1.5569738e-022 ub1=4.7964565e-020             lub1=-1.3595078e-025            wub1=-8.4388715e-025 pub1=1.8286553e-031             uc1=2.4672441e-010             luc1=9.5263544e-018 wuc1=2.9961842e-017             puc1=-3.0771844e-023            at=54626.485 lat=-0.0034176574              wat=0.011004466                pat=-2.1314863e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=2.0146756e-009             pkt2=-5.1331899e-030            lvsat=-0.0011956032 wvsat=0.0068219704               pvsat=-2.988023e-009             vth0_mcl=0.000194855 lvth0_mcl=-8.53466e-11               wvth0_mcl=-1.75623e-09               pvth0_mcl=7.69229e-16 vsat_ff=-7548.77                   vsat_ss=7757.96                    lvsat_ff=0.000678349 lvsat_ss=-0.000721022               wvsat_ff=-0.00175623                wvsat_ss=-0.000129141 pvsat_ff=7.69231e-10                pvsat_ss=-3.84611e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_12_mac.4 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=9.007e-06                  vth0=0.50515445 lvth0=-2.8978128e-009            wvth0=-2.3123211e-008            pvth0=2.6404181e-015 k2=-0.024410915               lk2=3.108119e-009              wk2=-1.5523557e-008 pk2=-6.8730342e-016            cit=0.00040041836              lcit=3.7097863e-010 wcit=1.3322287e-009             pcit=-1.8505113e-016            voff=-0.21716217 lvoff=-6.4778842e-010            wvoff=1.6658419e-008             pvoff=-2.7215737e-015 eta0=0.0094474074               weta0=-4.0293511e-009            etab=-0.050049327 wetab=4.4423596e-010             u0=0.02238272                 lu0=2.2734743e-010 wu0=-3.2103088e-010            pu0=-3.2867097e-017            ua=-1.4645625e-09 lua=3.4254463e-17              wua=-4.5406558e-17             pua=2.5913924e-24 ub=1.617192e-018              lub=-2.905358e-026             wub=3.35592e-026 pub=-1.5213525e-032            uc=4.6330271e-011             luc=7.2775811e-018 wuc=-2.2701853e-017            puc=-6.4007795e-024            vsat=90266.865 a0=2.9067412                  la0=-3.3918822e-007            wa0=-7.9388046e-007 pa0=1.0555337e-013             ags=-0.41052818                lags=2.7542615e-007 wags=1.5529311e-006             pags=-2.0582962e-013            keta=-0.07306067 lketa=-1.2071979e-008            wketa=-1.1032747e-008            pketa=6.3606185e-015 pclm=1.463455                   lpclm=6.3142857e-009             wpclm=5.0366889e-008 ppclm=3.0543433e-029             pdiblc2=0.007205798                lpdiblc2=-2.7109424e-010 wpdiblc2=3.6550637e-009             ppdiblc2=-2.4065038e-016            agidl=1.6334654e-010 lagidl=-3.5679975e-018            wagidl=-1.3996786e-017            pagidl=1.8379414e-025 aigbacc=0.013531                   aigc=0.011398772                laigc=-9.1083597e-012 waigc=2.7547407e-011             paigc=-5.2172465e-018            aigsd=0.010847082 laigsd=-1.9097642e-011            waigsd=1.4434095e-011             paigsd=3.5715255e-018 tvoff=0.00183399                 ltvoff=-8.97735e-012              wtvoff=-5.42144e-010 ptvoff=3.95711e-017               kt1=-0.16158242                lkt1=-2.1585121e-009 wkt1=-2.3626673e-008            pkt1=4.0950279e-015             kt2=-0.053401058 lkt2=-1.6781968e-010            ute=-0.47746913                lute=-4.0296298e-008 wute=-2.0905857e-007            pute=4.2647947e-014             ua1=1.8366289e-009 lua1=-1.5322215e-016            wua1=-1.7635027e-016            pua1=2.7009872e-023 ub1=-1.0865286e-018            lub1=9.5485817e-026             wub1=-6.9586414e-026 pub1=2.4908182e-032             uc1=3.9752127e-010             luc1=-2.1236206e-017 wuc1=-2.5557598e-016            puc1=2.7477872e-023             at=30541.866 lat=0.0014956049               wat=0.00092689141              pat=-7.5661008e-011 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=5.7562159e-009             pkt2=-7.6327422e-016            lvsat=0.0013468127 wvsat=-0.016666279               pvsat=1.8035799e-009             vth0_mcl=-0.000292692 lvth0_mcl=1.41131e-11                wvth0_mcl=2.63803e-09                pvth0_mcl=-1.27202e-16 vsat_ff=-6838.07                   vsat_ss=6838.07                    lvsat_ff=0.000533369 lvsat_ss=-0.000533369               wvsat_ff=0.00326157                 wvsat_ss=-0.00326157 pvsat_ff=-2.54402e-10               pvsat_ss=2.54402e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_12_mac.5 nmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=9e-007                     wmax=9.007e-06                  vth0=0.41703319 lvth0=3.9756459e-009             wvth0=1.2282915e-008             pvth0=-1.2125979e-016 k2=-0.010059655               lk2=1.9887206e-009             wk2=-2.3533657e-008 pk2=-6.2515596e-017            cit=0.0026372748               lcit=1.9650383e-010 wcit=-2.5284609e-009            pcit=1.1608266e-016             voff=-0.17613727 lvoff=-3.8477306e-009            wvoff=-2.919754e-008             pvoff=8.5519112e-016 eta0=0.0094474074               weta0=-4.0293511e-009            etab=-0.050049327 wetab=4.4423596e-010             u0=0.015244524                lu0=7.8412673e-010 wu0=8.3947763e-009             pu0=-7.1270006e-016            ua=-1.8635648e-09 lua=6.5376643e-17              wua=1.2082415e-16              pua=-1.0374602e-23 ub=1.3490388e-018             lub=-8.1376239e-027            wub=4.1996017e-025 pub=-4.53528e-032              uc=-5.7139095e-012            luc=1.1337027e-017 wuc=4.7456802e-017             puc=-1.1873155e-023            vsat=68093.215 a0=-1.5261505                 la0=6.5773376e-009             wa0=1.5468129e-006 pa0=-7.7020711e-014            ags=2.0756309                  lags=8.1505739e-008 wags=-3.6953403e-006            pags=2.0353555e-013             keta=-0.3810535 lketa=1.1951462e-008             wketa=8.9541136e-008             pketa=-1.4841443e-015 pclm=1.3555185                  lpclm=1.4733333e-008             wpclm=5.0366889e-008 ppclm=-2.2498332e-028            pdiblc2=0.0010072249               lpdiblc2=2.1239446e-010 wpdiblc2=-4.0495258e-009            ppdiblc2=3.603076e-016              agidl=9.0297202e-011 lagidl=2.1298511e-018             wagidl=-1.8923039e-017            pagidl=5.6804185e-025 aigbacc=0.013531                   aigc=0.011524806                laigc=-1.8938986e-011 waigc=-5.3884221e-011            paigc=1.1344206e-018             aigsd=0.010478405 laigsd=9.6591375e-012             waigsd=4.0761185e-011             paigsd=1.5180125e-018 tvoff=0.00181292                 ltvoff=-7.33423e-012              wtvoff=-6.76336e-010 ptvoff=5.0038e-017                kt1=-0.19197718                lkt1=2.1227932e-010 wkt1=3.7587059e-008             pkt1=-6.7964312e-016            kt2=-0.05470749 lkt2=-6.5918025e-011            ute=-1.1737326                 lute=1.4012251e-008 wute=5.9229782e-007             pute=-1.9857851e-014            ua1=7.8886156e-010 lua1=-7.1496297e-017            wua1=-3.3220617e-016            pua1=3.9166632e-023 ub1=-1.1252496e-018            lub1=9.8506056e-026             wub1=1.5307561e-024 pub1=-9.9918533e-032            uc1=-1.3520856e-010            luc1=2.0316721e-017 wuc1=4.0114429e-016             puc1=-2.3746309e-023            at=32617.669 lat=0.0013336923               wat=-0.00069448087             pat=5.080603e-011 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-1.1640348e-008            pkt2=5.9365773e-016             lvsat=0.0030763573 wvsat=0.0094805483               pvsat=-2.3587268e-010            vth0_mcl=-0.00241605 vth0_mc=-0.00314819                lvth0_mcl=1.79735e-10                lvth0_mc=2.45559e-10 wvth0_mcl=-3.74651e-09               wvth0_mc=2.85226e-09                pvth0_mcl=3.70794e-16 pvth0_mc=-2.22476e-16               u0_ff=0.000314272                u0_ss=-0.000125489 u0_mc=0.00209879                 lu0_ff=-2.45132e-11               lu0_ss=9.78822e-12 lu0_mc=-1.63706e-10               wu0_ff=5.70452e-10                wu0_ss=-5.70452e-10 wu0_mc=-1.90151e-09               pu0_ff=-4.44953e-17               pu0_ss=4.44952e-17 pu0_mc=1.48318e-16                vsat_ff=-210.974                   lvsat_ff=1.6456e-05 wvsat_ff=0.00190151                 pvsat_ff=-1.48318e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_12_mac.6 nmos ( level=54                         lmin=9e-007                     lmax=9.019e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=0.47766419 lvth0=2.3665305e-008             wvth0=-4.4574812e-009            pvth0=-8.1680085e-015 k2=-0.024493007               lk2=-8.3090004e-010            wk2=-4.3004223e-009 pk2=-1.1202063e-015            cit=0.003796706                lcit=-1.5093682e-009 wcit=-1.2554141e-009            pcit=1.0255895e-015             voff=-0.20186073 lvoff=-1.4960939e-008            wvoff=1.4126349e-009             pvoff=3.8182807e-015 eta0=0.0034833333               weta0=1.3741e-009                etab=-0.06140265 wetab=1.0730347e-008             u0=0.020131668                lu0=8.52511e-009 wu0=2.134362e-009              pu0=-5.2276819e-015            ua=-1.4217145e-009 lua=2.6579572e-016             wua=1.666244e-016              pua=-2.0148936e-022 ub=1.7957089e-018             lub=2.4755469e-025             wub=-3.0759686e-026 pub=-1.6938177e-031            uc=9.4602594e-011             luc=5.0682735e-017 wuc=-1.7045601e-018            puc=-3.8669821e-023            vsat=100000 a0=1.2680021                  la0=1.0392934e-006             wa0=6.8592501e-008 pa0=-2.7763191e-013            ags=0.4635759                  lags=8.8967675e-007 wags=5.5472982e-008             pags=-2.5527877e-013            keta=0.0071807891 lketa=-6.4540933e-008            wketa=-2.1623886e-009            pketa=1.9435549e-014 pclm=1.1837383                  lpclm=1.4616041e-007             wpclm=-1.5064207e-008 ppclm=1.353971e-013              pdiblc2=0.0010234936               lpdiblc2=2.8771024e-009 wpdiblc2=-1.3978198e-010            ppdiblc2=9.4399604e-016             agidl=1.7682491e-010 lagidl=-2.0044097e-017            wagidl=-2.280406e-017             pagidl=1.3773386e-023 aigbacc=0.013531                   aigc=0.011448965                laigc=-6.6368636e-011 waigc=-1.8500835e-011            paigc=2.1367016e-017             aigsd=0.010825399 laigsd=1.084341e-010              waigsd=1.2591647e-011             paigsd=-5.5400971e-017 tvoff=0.00177287                 ltvoff=2.36057e-010               wtvoff=1.88392e-011 ptvoff=-2.82829e-016              kt1=-0.14099914                lkt1=7.2113404e-009 wkt1=-3.3521742e-009            pkt1=-1.1376931e-014            kt2=-0.067886716 lkt2=-1.0181961e-009            ute=-1.0308146                 lute=2.649128e-007 wute=2.2047756e-007             pute=-1.6947654e-013            ua1=9.3466812e-010 lua1=4.7450718e-016             wua1=5.3390012e-016             pua1=-4.5189616e-022 ub1=-6.8553279e-019            lub1=2.9095316e-025             wub1=-9.0375616e-026 pub1=-1.388091e-031             uc1=2.049843e-010              luc1=2.7038034e-016 wuc1=9.8642059e-017             puc1=-1.9497182e-022            at=123288.06 lat=-0.029553044               wat=-0.001434336               pat=1.2891812e-008 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-3.0128415e-010            pkt2=2.7079419e-015             lvsat=0 wvsat=0                          pvsat=0                          ags_ff=0.133495 ags_ss=-0.116669                  ags_fs=0.0944821                  ags_sf=-0.100213 lags_ff=-1.18543e-07               lags_ss=1.03602e-07                lags_fs=-8.38998e-08 lags_sf=8.89899e-08                wags_ff=-3.04877e-08               wags_ss=1.52438e-08 wags_fs=-1.52436e-08               wags_sf=3.04878e-08                pags_ff=2.70729e-14 pags_ss=-1.35364e-14               pags_fs=1.35366e-14                pags_sf=-2.70732e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.7 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.51001587 lvth0=-5.0629897e-009            wvth0=-2.1283387e-008            pvth0=6.7733962e-015 k2=-0.023728576               lk2=-1.5097146e-009            wk2=-6.3647135e-009 pk2=7.1288432e-016             cit=0.0011679689               lcit=8.2495035e-010 wcit=4.1705274e-010             pcit=-4.5956098e-016            voff=-0.21707295 lvoff=-1.4524864e-009            wvoff=9.3869453e-009             pvoff=-3.2629069e-015 eta0=0.0034833333               weta0=1.3741e-009                etab=-0.06140265 wetab=1.0730347e-008             u0=0.03318417                 lu0=-3.0655126e-009 wu0=-5.8979487e-009            pu0=1.90501e-015               ua=-1.0179958e-009 lua=-9.2706409e-017            wua=-7.3328978e-017            pua=1.1589243e-023 ub=2.3507349e-018             lub=-2.4530842e-025            wub=-3.5123828e-025 pub=1.1520323e-031             uc=2.2690859e-010             luc=-6.6804986e-017 wuc=-8.0948973e-017            puc=3.1699218e-023             vsat=100000 a0=3.0502815                  la0=-5.4337075e-007            wa0=-6.3145424e-007 pa0=3.440096e-013              ags=1.7084002                  lags=-2.1572721e-007 wags=-5.7538991e-007            pags=3.0492747e-013             keta=-0.067502288 lketa=1.7776394e-009             wketa=3.8421449e-008             pketa=-1.6602899e-014 pclm=1.3483333                  lpclm=0                          wpclm=1.3741e-007 ppclm=0                          pdiblc2=0.0053264193               lpdiblc2=-9.4389554e-010 wpdiblc2=6.3894108e-010             ppdiblc2=2.5248997e-016             agidl=1.5136405e-010 lagidl=2.5651399e-018             wagidl=3.4481308e-018             pagidl=-9.5385598e-024 aigbacc=0.013531                   aigc=0.011380727                laigc=-5.7732917e-012 waigc=2.7189678e-011             paigc=-1.9206159e-017            aigsd=0.011170278 laigsd=-1.9781778e-010            waigsd=-1.3310558e-010            paigsd=7.3978167e-017 tvoff=0.00258686                 ltvoff=-4.86762e-010              wtvoff=-6.15026e-010 ptvoff=2.80043e-016               kt1=-0.097338048               lkt1=-3.1559707e-008 wkt1=-3.4737673e-008            pkt1=1.6493393e-014             kt2=-0.090511556 lkt2=1.9072661e-008             ute=-0.69230056                lute=-3.5687629e-008 wute=5.9659758e-009             pute=2.1009743e-014             ua1=1.2301045e-009 lua1=2.1215963e-016             wua1=3.3999245e-016             pua1=-2.7970615e-022 ub1=4.5912197e-019             lub1=-7.2550027e-025            wub1=-8.9617483e-025 pub1=5.767406e-031              uc1=8.1094044e-010             luc1=-2.6770871e-016 wuc1=-2.6001636e-016            puc1=1.2351686e-022             at=109033.04 lat=-0.016894594               wat=0.040687984                pat=-2.4512809e-008 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=8.0980293e-009             pkt2=-4.7506485e-015            lvsat=0 wvsat=0                          pvsat=0                          vsat_ff=7316.19 vsat_ss=-9295.36                   lvsat_ff=-0.00649677                lvsat_ss=0.00825423 wvsat_ff=-0.00133745                wvsat_ss=0.00401238                 pvsat_ff=1.18766e-09 pvsat_ss=-3.56299e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.8 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.51110662 lvth0=-5.5407385e-009            wvth0=-7.5487085e-009            pvth0=7.5760682e-016 k2=-0.026944473               lk2=-1.0115215e-010            wk2=-6.8231326e-009 pk2=9.1367189e-016             cit=0.0032658385               lcit=-9.3916556e-011 wcit=-1.0906496e-009            pcit=2.0081266e-016             voff=-0.22918309 lvoff=3.8517574e-009             wvoff=8.6609619e-009             pvoff=-2.9449262e-015 eta0=0.0034833333               weta0=1.3741e-009                etab=-0.062216891 wetab=1.1468049e-008             u0=0.026744932                lu0=-2.4512614e-010 wu0=-8.621949e-010             pu0=-3.0065012e-016            ua=-1.281528e-009 lua=2.2720677e-017             wua=4.0693429e-017             pua=-3.8352572e-023 ub=2.1061973e-018             lub=-1.3820094e-025            wub=-1.6572351e-025 pub=3.3947754e-032             uc=1.31296e-010               luc=-2.4926675e-017 wuc=-2.6486427e-017            puc=7.8446228e-024             vsat=121324.08 a0=2.8427095                  la0=-4.524542e-007             wa0=4.0073958e-008 pa0=4.9880247e-014             ags=0.21929943                 lags=4.3649892e-007 wags=8.7298098e-007             pags=-3.2945898e-013            keta=-0.0063284722 lketa=-2.5016492e-008            wketa=-1.4009654e-008            pketa=6.3619245e-015 pclm=1.1725214                  lpclm=7.7005641e-008             wpclm=2.5720333e-007 ppclm=-5.246948e-014             pdiblc2=-0.0011399712              lpdiblc2=1.8883835e-009 wpdiblc2=1.8861194e-009             ppdiblc2=-2.9377412e-016            agidl=1.7520875e-010 lagidl=-7.878839e-018             wagidl=-3.0213374e-017            pagidl=5.2051791e-024 aigbacc=0.013531                   aigc=0.011337219                laigc=1.3283507e-011 waigc=5.1752094e-012             paigc=-9.563822e-018             aigsd=0.010743129 laigsd=-1.0726741e-011            waigsd=-1.0543156e-011            paigsd=2.0295825e-017 tvoff=0.00121119                 ltvoff=1.1578e-010                wtvoff=3.40221e-010 ptvoff=-1.38355e-016              kt1=-0.17283151                lkt1=1.5064299e-009 wkt1=1.3865128e-008             pkt1=-4.7946343e-015            kt2=-0.039934188 lkt2=-3.0802256e-009            ute=-0.92751278                lute=6.7335323e-008 wute=1.6221462e-007             pute=-4.7427163e-014            ua1=2.3516441e-009 lua1=-2.790747e-016             wua1=-6.0110733e-016            pua1=1.3249555e-022 ub1=-2.0495219e-018            lub1=3.7328574e-025             wub1=1.0564356e-024 pub1=-2.7850275e-031            uc1=1.7090598e-010             luc1=1.2626379e-017 wuc1=9.8653333e-017             puc1=-3.3580467e-023            at=101356.94 lat=-0.013532462               wat=-0.031333329               pat=7.0325266e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-7.5399333e-009            pkt2=2.0987792e-015             lvsat=-0.0093399455 wvsat=-0.010024546               pvsat=4.390751e-009              letab=3.5663755e-010 petab=-3.2311362e-016            vth0_mcl=-0.00174359                lvth0_mcl=7.63693e-10 wvth0_mcl=3.3e-15                    pvth0_mcl=-4e-22                     vsat_ff=-13648.3 vsat_ss=16132                      lvsat_ff=0.00268565                 lvsat_ss=-0.00288294 wvsat_ff=0.00376993                 wvsat_ss=-0.0077161                 pvsat_ff=-1.04939e-09 pvsat_ss=1.57408e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.9 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.48463779 lvth0=-1.4109765e-010            wvth0=-4.5351169e-009            pvth0=1.4283414e-016 k2=-0.042591293               lk2=3.0907993e-009             wk2=9.4786576e-010 pk2=-6.7161178e-016            cit=0.0026656504               lcit=2.8521826e-011 wcit=-7.2007156e-010            pcit=1.2521473e-016             voff=-0.19044289 lvoff=-4.0512431e-009            wvoff=-7.5492459e-009            pvoff=3.6195623e-016 eta0=0.0034833333               weta0=1.3741e-009                etab=-0.059890488 wetab=9.3603283e-009             u0=0.023186175                lu0=4.8086022e-010 wu0=-1.0489618e-009            pu0=-2.6254968e-016            ua=-1.2965046e-09 lua=2.5775891e-17              wua=-1.9766711e-16             pua=1.0272979e-23 ub=1.4787573e-018             lub=-1.0203183e-026            wub=1.5898109e-025 pub=-3.2291985e-032            uc=-1.2983305e-011            luc=4.5063042e-018 wuc=3.1036246e-017             puc=-3.8900027e-024            vsat=54670.318 a0=1.1223615                  la0=-1.0150321e-007            wa0=8.2276756e-007 pa0=-1.0978925e-013            ags=3.1722016                  lags=-1.6589312e-007 wags=-1.6930221e-006            pags=1.9400565e-013             keta=-0.12532143 lketa=-7.4192857e-010            wketa=3.63155e-008               pketa=-3.904407e-015 pclm=1.4251587                  lpclm=2.5467619e-008             wpclm=8.5063333e-008 ppclm=-1.735292e-014             pdiblc2=0.0089603323               lpdiblc2=-1.7207842e-010 wpdiblc2=2.0654556e-009             ppdiblc2=-3.3035871e-016            agidl=1.6232592e-010 lagidl=-5.2507411e-018            wagidl=-1.3072103e-017            pagidl=1.7083599e-024 aigbacc=0.013531                   aigc=0.011491412                laigc=-1.8171894e-011 waigc=-5.6384289e-011            paigc=2.9943158e-018             aigsd=0.010675017 laigsd=3.1681838e-012             waigsd=1.7032516e-010             paigsd=-1.6601313e-017 tvoff=0.00160732                 ltvoff=3.49699e-011               wtvoff=-3.36787e-010 ptvoff=-2.45157e-019              kt1=-0.19543154                lkt1=6.1168359e-009 wkt1=7.0406331e-009             pkt1=-3.4024374e-015            kt2=-0.048203175 lkt2=-1.3933524e-009            ute=-0.63302176                lute=7.2591554e-009 wute=-6.8127878e-008            pute=-4.3729358e-016            ua1=1.6881169e-009 lua1=-1.4371515e-016            wua1=-4.1798381e-017            pua1=1.8396527e-023 ub1=-8.5044715e-019            lub1=1.2867449e-025             wub1=-2.8347618e-025 pub1=-5.1607584e-033            uc1=1.5818413e-010             luc1=1.5221638e-017 wuc1=-3.8736533e-017            puc1=-5.5529344e-024            at=30165.477 lat=0.00099059728              wat=0.0012678999               pat=3.8187589e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=1.0469333e-009             pkt2=3.470584e-016              lvsat=0.0042574213 wvsat=0.015584193                pvsat=-8.334316e-010             letab=-1.1794862e-010 petab=1.0686145e-016             vth0_mcl=0.00261905                 lvth0_mcl=-1.26285e-10 wvth0_mcl=-3.33e-15                  pvth0_mcl=-8e-22                     vsat_ff=-782.543 vsat_ss=3238.1                     lvsat_ff=6.1038e-05                 lvsat_ss=-0.000252571 wvsat_ff=-0.00222473                wvsat_ss=-3.3e-09                   pvsat_ff=1.7353e-10 pvsat_ss=-4e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.10 nmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.414403 lvth0=5.3372164e-009             wvth0=1.4665867e-008             pvth0=-1.3548426e-015 k2=-0.028547711               lk2=1.9953999e-009             wk2=-6.783478e-009 pk2=-6.8566966e-017            cit=-0.0026574729              lcit=4.4372544e-010 wcit=2.2685805e-009             pcit=-1.0790012e-016            voff=-0.19709715 lvoff=-3.5322108e-009            wvoff=-1.0207886e-008            pvoff=5.6933013e-016 eta0=0.0034833333               weta0=1.3741e-009                etab=-0.06140265 wetab=1.0730347e-008             u0=0.03291506                 lu0=-2.7799282e-010 wu0=-7.6147301e-009            pu0=2.4958025e-016             ua=-1.8481297e-09 lua=6.8802645e-17              wua=1.068398e-16               pua=-1.3478561e-23 ub=2.6777321e-018             lub=-1.0372322e-025            wub=-7.8383598e-025 pub=4.1247747e-032             uc=5.5445981e-011             luc=-8.3118003e-019 wuc=-7.9540589e-018            puc=-8.4875889e-025            vsat=53583.632 a0=-1.8819064                 la0=1.3282969e-007             wa0=1.8691277e-006 pa0=-1.9140534e-013            ags=-4.5356074                 lags=4.3531598e-007 wags=2.2944416e-006             pags=-1.1701652e-013            keta=-0.353 lketa=1.7017e-008                wketa=6.4124667e-008             pketa=-6.073522e-015 pclm=1.8492593                  lpclm=-7.6122222e-009            wpclm=-3.9696222e-007 ppclm=2.0245073e-014             pdiblc2=-0.00084064828             lpdiblc2=5.9239806e-010 wpdiblc2=-2.3753527e-009            ppdiblc2=1.6024338e-017             agidl=2.6028575e-011 lagidl=5.3804518e-018             wagidl=3.9304337e-017             pagidl=-2.3770024e-024 aigbacc=0.013531                   aigc=0.011529478                laigc=-2.1141042e-011 waigc=-5.8117208e-011            paigc=3.1294834e-018             aigsd=0.010635792 laigsd=6.22775e-012               waigsd=-1.0183077e-010            paigsd=4.6268496e-018 tvoff=0.000903737                ltvoff=8.98496e-011               wtvoff=1.47384e-010 ptvoff=-3.80105e-017              kt1=-0.10476229                lkt1=-9.5536557e-010 wkt1=-4.142963e-008             pkt1=3.7824316e-016             kt2=-0.085081482 lkt2=1.4831556e-009             ute=-0.98898611                lute=3.5024375e-008 wute=4.2491752e-007             pute=-3.8894835e-014            ua1=-2.7376289e-010 lua1=9.3114755e-018             wua1=6.3053158e-016             pua1=-3.404521e-023 ub1=9.7495439e-019             lub1=-1.3706828e-026            wub1=-3.7202872e-025 pub1=1.74634e-033               uc1=4.9764444e-010             luc1=-1.1256267e-017 wuc1=-1.7222053e-016            puc1=4.8588176e-024             at=14112.377 lat=0.0022427391               wat=0.016071313                pat=-7.7279036e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=1.5878489e-008             pkt2=-8.0980293e-016            lvsat=0.0043421828 wvsat=0.022626231                pvsat=-1.3827106e-009            vth0_mcl=-0.000824851 lvth0_mcl=1.42337e-10                wvth0_mcl=-5.18807e-09               pvth0_mcl=4.04673e-16 cit_mcl=0.000286319                lcit_mcl=-2.23329e-11               wcit_mcl=-2.59405e-10 pcit_mcl=2.02336e-17                voff_mcl=-0.00286319                lvoff_mcl=2.23329e-10 wvoff_mcl=2.59405e-09                pvoff_mcl=-2.02336e-16               u0_ss=-0.000755123 u0_ff=0.000800754                lu0_ss=5.89004e-11                lu0_ff=-6.2458e-11 wu0_ss=-1e-15                     wu0_ff=1.29699e-10                pu0_ss=3.9e-23 pu0_ff=-1.01169e-17               vsat_ff=10477.4                    vsat_fs=2863.19 vsat_ss=2863.19                    lvsat_ff=-0.000817237               lvsat_fs=-0.000223329 lvsat_ss=-0.000223329               wvsat_ff=-0.00778216                wvsat_fs=-0.00259405 wvsat_ss=-0.00259405                pvsat_ff=6.07008e-10                pvsat_fs=2.02336e-10 pvsat_ss=2.02336e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.11 nmos ( level=54                         lmin=9e-007                     lmax=9.019e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.47341668 lvth0=7.4321438e-009             wvth0=-2.1383439e-009            pvth0=6.9529727e-016 k2=-0.031842039               lk2=-1.1526374e-009            wk2=-2.8785119e-010 pk2=-9.4453764e-016            cit=0.0013365725               lcit=9.0110111e-010 wcit=8.7818848e-011             pcit=-2.9052672e-016            voff=-0.20846642 lvoff=-5.2653687e-009            wvoff=5.0193458e-009             pvoff=-1.4755008e-015 eta0=0.0039555556               weta0=1.1162667e-009             etab=-0.044893333 wetab=1.71626e-009               u0=0.025279907                lu0=-3.6239243e-009 wu0=-6.7657667e-010            pu0=1.4056909e-015             ua=-1.0485726e-009 lua=-2.1287643e-016            wua=-3.7111016e-017            pua=5.9865629e-023 ub=1.7329505e-018             lub=-5.823644e-026             wub=3.5064003e-027 pub=-2.4198121e-033            uc=8.9513149e-011             luc=-2.6756617e-017 wuc=1.0742769e-018             puc=3.6120652e-024             vsat=104088.89 a0=1.4442137                  la0=4.3111767e-007             wa0=-2.7619013e-008 pa0=5.4432035e-014             ags=0.56253859                 lags=2.1742994e-007 wags=1.4393494e-009             pags=1.1176798e-013             keta=0.012091527 lketa=-1.6801309e-008            wketa=-4.8436514e-009            pketa=-6.6302852e-015 pclm=1.133735                   lpclm=5.9559001e-007             wpclm=1.223759e-008 ppclm=-1.0999146e-013            pdiblc2=0.0010856629               lpdiblc2=2.820775e-009 wpdiblc2=-1.7372642e-010            ppdiblc2=9.7475084e-016             agidl=1.3393939e-010 lagidl=5.8487139e-018             wagidl=6.1142849e-019             pagidl=-3.6408878e-025 aigbacc=0.013531                   aigc=0.011442978                laigc=-1.8049513e-011 waigc=-1.5231601e-011            paigc=-5.0152256e-018            aigsd=0.010845286 laigsd=5.0945374e-011             waigsd=1.7337446e-012             paigsd=-2.4012126e-017 tvoff=0.00183037                 ltvoff=-4.67646e-010              wtvoff=-1.25558e-011 ptvoff=1.01393e-016               kt1=-0.14793959                lkt1=-1.0832969e-008 wkt1=4.3731104e-010             pkt1=-1.5247374e-015            kt2=-0.070482963 lkt2=3.9414044e-009             ute=-0.6010353                 lute=-7.1480873e-008 wute=-1.4181912e-008            pute=1.4194398e-014             ua1=2.102001e-009 lua1=-5.714233e-016             wua1=-1.0346366e-016            pua1=1.1918188e-022 ub1=-9.0317819e-019            lub1=8.4860408e-026             wub1=2.8458772e-026 pub1=-2.6282459e-032            uc1=4.3919671e-010             luc1=-1.2700081e-016 wuc1=-2.9237918e-017            puc1=2.1998292e-023             at=120172.9 lat=-0.0015540555              wat=0.00026653716              pat=-2.395636e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=1.1162667e-009             pkt2=-6.8207409e-030            lvsat=0 wvsat=-0.0022325333              pvsat=0                          ags_ff=0.0889965 ags_ss=-0.0774097                 ags_fs=0.134604                   ags_sf=-0.0216945 lags_ff=-7.90291e-08               lags_ss=6.87397e-08                lags_fs=-1.19528e-07 lags_sf=1.92646e-08                wags_ff=-6.19181e-09               wags_ss=-6.19183e-09 wags_fs=-3.71507e-08               wags_sf=-1.23836e-08               pags_ff=5.49829e-15 pags_ss=5.49831e-15                pags_fs=3.29898e-14                pags_sf=1.09966e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.12 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.46989219 lvth0=1.0561894e-008             wvth0=6.2414209e-010             pvth0=-1.7577903e-015 k2=-0.032370158               lk2=-6.8366736e-010            wk2=-1.6464099e-009 pk2=2.6186251e-016             cit=0.0028528431               lcit=-4.4534716e-010 wcit=-5.0288856e-010            pcit=2.3402146e-016             voff=-0.20130231 lvoff=-1.1627102e-008            wvoff=7.7617664e-010             pvoff=2.2924334e-015 eta0=0.0039555556               weta0=1.1162667e-009             etab=-0.044893333 wetab=1.71626e-009               u0=0.019853658                lu0=1.1945851e-009 wu0=1.3805113e-009             pu0=-4.2100326e-016            ua=-1.2778753e-009 lua=-9.2556781e-018            wua=6.8565207e-017             pua=-3.3974857e-023 ub=1.7245165e-018             lub=-5.0747108e-026            wub=-9.3230592e-027 pub=8.9727479e-033             uc=6.6249583e-011             luc=-6.0985704e-018 wuc=6.7708421e-018             puc=-1.4464847e-024            vsat=104088.89 a0=1.6353582                  la0=2.6138129e-007             wa0=1.4109388e-007 pa0=-9.5385019e-014            ags=0.38245718                 lags=3.7734224e-007 wags=1.4857497e-007             pags=-1.8888445e-014            keta=0.039895481 lketa=-4.1491221e-008            wketa=-2.0217733e-008            pketa=7.0218989e-015 pclm=1.9039407                  lpclm=-8.8352711e-008            wpclm=-1.6595164e-007 ppclm=4.824058e-014              pdiblc2=0.0049111762               lpdiblc2=-5.7628081e-010 wpdiblc2=8.6566379e-010             ppdiblc2=5.1772326e-017             agidl=1.6423652e-010 lagidl=-2.105513e-017             wagidl=-3.5802344e-018            pagidl=3.3581078e-024 aigbacc=0.013531                   aigc=0.011486035                laigc=-5.6284434e-011 waigc=-3.0308346e-011            paigc=8.3729246e-018             aigsd=0.011024483 laigsd=-1.0818178e-010            waigsd=-5.3501655e-011            paigsd=2.5036909e-017 tvoff=0.00126551                 ltvoff=3.39546e-011               wtvoff=1.06432e-010 ptvoff=-4.2677e-018               kt1=-0.15282388                lkt1=-6.4957136e-009 wkt1=-4.442407e-009             pkt1=2.8084522e-015             kt2=-0.07971437 lkt2=1.2138894e-008             ute=-0.68788938                lute=5.6455462e-009 wute=3.5574674e-009             pute=-1.5581707e-015            ua1=1.7289049e-009 lua1=-2.401139e-016             wua1=6.7647469e-017             pua1=-3.2764799e-023 ub1=-1.1882276e-018            lub1=3.3798427e-025             wub1=3.2780287e-027 pub1=-3.9219592e-033            uc1=3.5085748e-010             luc1=-4.8555577e-017 wuc1=-8.8110649e-018            puc1=3.8592464e-024             at=197133.1 lat=-0.069894709               wat=-0.0074146454              pat=4.4252541e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=2.2027662e-009             pkt2=-9.6481161e-016            lvsat=0 wvsat=-0.0022325333              pvsat=0                          vsat_ff=9841.48 vsat_ss=-3936.59                   lvsat_ff=-0.00873924                lvsat_ss=0.00349569 wvsat_ff=-0.00271625                wvsat_ss=0.0010865                  pvsat_ff=2.41203e-09 pvsat_ss=-9.64812e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.13 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.51389535 lvth0=-8.7114913e-009            wvth0=-9.0713559e-009            pvth0=2.4888378e-015 k2=-0.038205269               lk2=1.872111e-009              wk2=-6.7473804e-010 pk2=-1.6372977e-016            cit=0.00077646505              lcit=4.6410641e-010 wcit=2.6854827e-010             pcit=-1.0386788e-016            voff=-0.23086584 lvoff=1.3217237e-009             wvoff=9.5797409e-009             pvoff=-1.5635277e-015 eta0=0.0039555556               weta0=1.1162667e-009             etab=-0.043807679 wetab=1.4166193e-009             u0=0.024084788                lu0=-6.5865013e-010 wu0=5.9024363e-010             pu0=-7.4866021e-017            ua=-1.2577297e-009 lua=-1.8079465e-017            wua=2.769954e-017              pua=-1.6075694e-023 ub=1.8514737e-018             lub=-1.0635434e-025            wub=-2.6644427e-026 pub=1.6559507e-032             uc=6.9001586e-011             luc=-7.3039478e-018 wuc=7.5263247e-018             puc=-1.7773861e-024            vsat=111622.9 a0=2.7811947                  la0=-2.404951e-007             wa0=7.3661016e-008 pa0=-6.5849422e-014            ags=1.9022442                  lags=-2.8832449e-007 wags=-4.5906876e-008            pags=6.6294603e-014             keta=-0.037688034 lketa=-7.509641e-009             wketa=3.1126667e-009             pketa=-3.196816e-015 pclm=1.8349288                  lpclm=-5.812547e-008             wpclm=-1.0447111e-007 ppclm=2.1312107e-014             pdiblc2=0.0008417676               lpdiblc2=1.2061202e-009 wpdiblc2=8.0408996e-010             ppdiblc2=7.8741666e-017             agidl=1.0706074e-010 lagidl=3.9878605e-018             wagidl=6.9954429e-018             pagidl=-1.2740388e-024 aigbacc=0.013531                   aigc=0.01135168                 laigc=2.5631796e-012 waigc=-2.7205665e-012            paigc=-3.710523e-018             aigsd=0.010651841 laigsd=5.5035485e-011             waigsd=3.9300309e-011             paigsd=-1.5610351e-017 tvoff=0.00166224                 ltvoff=-1.39814e-010              wtvoff=9.39501e-011 ptvoff=1.19938e-018               kt1=-0.16087903                lkt1=-2.9675578e-009 wkt1=7.3390753e-009             pkt1=-2.351837e-015             kt2=-0.055525926 lkt2=1.5443556e-009             ute=-0.6437572                 lute=-1.3684348e-008 wute=7.2840693e-009             pute=-3.1904224e-015            ua1=1.1662854e-009 lua1=6.3134484e-018             wua1=4.6098551e-017             pua1=-2.3326373e-023 ub1=2.4939345e-020             lub1=-1.9338285e-025            wub1=-7.6220262e-026 pub1=3.0898292e-032             uc1=3.5871909e-010             luc1=-5.1998961e-017 wuc1=-3.8926222e-018            puc1=1.7049685e-024             at=40570.026 lat=-0.0013200829              wat=0.0018563282               pat=3.6456767e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=9.7315556e-010             pkt2=-4.2624213e-016            lvsat=-0.0032998975 wvsat=-0.0047277042              pvsat=1.0928848e-009             letab=-4.7551673e-010 petab=1.3124262e-016             vth0_mcl=-0.00263476                lvth0_mcl=1.15403e-09 wvth0_mcl=4.86578e-10                pvth0_mcl=-2.13121e-16               vsat_ff=-14082.6 vsat_ss=4044.44                    lvsat_ff=0.00173953                 lvsat_ss=-4.4e-09 wvsat_ff=0.00400712                 wvsat_ss=-0.00111626                pvsat_ff=-5.32808e-10 pvsat_ss=-1.3e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.14 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.47311032 lvth0=-3.9134488e-010            wvth0=1.7588829e-009             pvth0=2.7946913e-016 k2=-0.038159319               lk2=1.8627373e-009             wk2=-1.4719923e-009 pk2=-1.0899053e-018            cit=0.0019221001               lcit=2.3039685e-010 wcit=-3.1409312e-010            pcit=1.4990967e-017             voff=-0.20836025 lvoff=-3.2694166e-009            wvoff=2.2336294e-009             pvoff=-6.4921014e-017 eta0=0.0039555556               weta0=1.1162667e-009             etab=-0.046909549 wetab=2.2727355e-009             u0=0.022067931                lu0=-2.472113e-010 wu0=-4.3840044e-010            pu0=1.3497737e-016             ua=-1.5833178e-09 lua=4.8340496e-17              wua=-4.1067123e-17             pua=-2.0472952e-24 ub=1.7730302e-018             lub=-9.0351872e-026            wub=-1.6919413e-027 pub=1.14692e-032               uc=5.0989294e-011             luc=-3.6294403e-018 wuc=-3.8927925e-018            puc=5.5211381e-025             vsat=84818.008 a0=3.3537839                  la0=-3.573033e-007             wa0=-3.9558909e-007 pa0=2.9877599e-014             ags=-1.0724868                 lags=3.1852063e-007 wags=6.2457778e-007             pags=-7.0484267e-014            keta=-0.034227513 lketa=-8.2155873e-009            wketa=-1.3421778e-008            pketa=1.7621067e-016 pclm=1.6125926                  lpclm=-1.2768889e-008            wpclm=-1.7275556e-008 ppclm=3.5242133e-015             pdiblc2=0.0085545932               lpdiblc2=-3.6729627e-010 wpdiblc2=2.2869891e-009             ppdiblc2=-2.2376976e-016            agidl=1.3988975e-010 lagidl=-2.7092572e-018            wagidl=-8.2195166e-019            pagidl=3.2070969e-025 aigbacc=0.013531                   aigc=0.011436407                laigc=-1.472118e-011 waigc=-2.6351689e-011            paigc=1.1102259e-018             aigsd=0.01112901 laigsd=-4.2306997e-011            waigsd=-7.7555019e-011            paigsd=8.2281359e-018 tvoff=0.000770921                ltvoff=4.20155e-011               wtvoff=1.19888e-010 ptvoff=-4.09204e-018              kt1=-0.16896492                lkt1=-1.3180376e-009 wkt1=-7.4101433e-009            pkt1=6.5700359e-016             kt2=-0.04424127 lkt2=-7.5771429e-010            ute=-0.73302235                lute=4.5257432e-009 wute=-1.3527557e-008            pute=1.0551495e-015             ua1=1.7499826e-009 lua1=-1.1276079e-016            wua1=-7.5577036e-017            pua1=1.4954462e-024 ub1=-1.4871713e-018            lub1=1.1508774e-025             wub1=6.4175234e-026 pub1=2.2576111e-033             uc1=9.8044444e-011             luc1=1.1786667e-018 wuc1=-5.9002667e-018            puc1=2.114528e-024              at=23452.328 lat=0.0021719274               wat=0.0049332792               pat=-2.6313033e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-1.1162667e-009            pkt2=1.1031247e-030             lvsat=0.0021683007 wvsat=-0.00087644634             pvsat=3.0722823e-010             letab=1.5726483e-010 petab=-4.3405093e-017            vth0_mcl=0.00427407                 lvth0_mcl=-2.55378e-10 wvth0_mcl=-9.03646e-10               pvth0_mcl=7.04847e-17                vsat_ff=-8994.71 vsat_ss=6548.15                    lvsat_ff=0.000701587                lvsat_ss=-0.000510756 wvsat_ff=0.00225911                 wvsat_ss=-0.00180729                pvsat_ff=-1.76211e-10 pvsat_ss=1.40969e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.15 nmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.43661491 lvth0=2.4552974e-009             wvth0=2.5381652e-009             pvth0=2.1868511e-016 k2=-0.040012067               lk2=2.0072516e-009             wk2=-5.2393959e-010 pk2=-7.5038015e-017            cit=0.0011727432               lcit=2.888467e-010 wcit=1.7728251e-010             pcit=-2.3336332e-017            voff=-0.23255497 lvoff=-1.3822287e-009            wvoff=9.1520787e-009             pvoff=-6.0456006e-016 eta0=0.0039555556               weta0=1.1162667e-009             etab=-0.044893167 wetab=1.716169e-009              u0=0.016513974                lu0=1.8599738e-010 wu0=1.3402632e-009             pu0=-3.7583973e-018            ua=-1.507223e-09 lua=4.240511e-17               wua=-7.929518e-17              pua=9.3449325e-25 ub=8.846418e-019              lub=-2.1057575e-026            wub=1.951913e-025 pub=-3.8876932e-033            uc=6.6309062e-011             luc=-4.8243822e-018 wuc=-1.3885301e-017            puc=1.3315295e-024             vsat=108541.49 a0=5.909353                   la0=-5.5663768e-007            wa0=-2.3848999e-006 pa0=1.8504384e-013             ags=-0.094280988               lags=2.4222058e-007 wags=-1.3052258e-007            pags=-1.1586439e-014            keta=-0.099259259 lketa=-3.1431111e-009            wketa=-7.4417778e-008            pketa=4.9338987e-015 pclm=0.9745679                  lpclm=3.6997037e-008             wpclm=8.0619259e-008 ppclm=-4.1115822e-015            pdiblc2=-0.0070620764              lpdiblc2=8.5080396e-010 wpdiblc2=1.021547e-009              ppdiblc2=-1.2506528e-016            agidl=9.912805e-011 lagidl=4.701551e-019              wagidl=-6.0797619e-019            pagidl=3.040196e-025 aigbacc=0.0055885832               aigc=0.011437817                laigc=-1.4831175e-011 waigc=-8.0705398e-012            paigc=-3.1570373e-019            aigsd=0.01035543 laigsd=1.803226e-011              waigsd=5.1246891e-011             paigsd=-1.818413e-018 tvoff=0.00134151                 ltvoff=-2.49085e-012              wtvoff=-9.16428e-011 ptvoff=1.24074e-017               kt1=-0.11109489                lkt1=-5.8318995e-009 wkt1=-3.7972029e-008            pkt1=3.0408307e-015             kt2=-0.053955556 ute=0.42525847                 lute=-8.5820161e-008            wute=-3.4726002e-007 pute=2.7086281e-014             ua1=1.2435061e-009             lua1=-7.3255624e-017 wua1=-1.978973e-016             pua1=1.1036427e-023             ub1=5.6046125e-019 lub1=-4.4627607e-026            wub1=-1.4571547e-025            pub1=1.8629086e-032 uc1=2.7081481e-010             luc1=-1.2297422e-017            wuc1=-4.8371556e-017 puc1=5.4272885e-024             at=32215.115                  lat=0.00148843 wat=0.0061872186               pat=-3.609376e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-1.1162667e-009            lvsat=0.0003178691               wvsat=-0.0073807602 pvsat=8.1456471e-010             letab=-1.2997419e-014            petab=7.0965909e-021 laigbacc=6.1950851e-010             waigbacc=4.3365596e-009             paigbacc=-3.3825165e-016 vth0_mcl=-0.018046                  lvth0_mcl=1.48558e-09                wvth0_mcl=4.21462e-09 pvth0_mcl=-3.28741e-16               cit_mcl=0.000390149                lcit_mcl=-3.04317e-11 wcit_mcl=-3.16097e-10               pcit_mcl=2.46555e-17                voff_mcl=-4.19517e-05 lvoff_mcl=3.27226e-12                wvoff_mcl=1.05366e-09                pvoff_mcl=-8.21851e-17 u0_ff=0.000941808                u0_ss=-0.000369178               u0_mc=-0.00154382 lu0_ff=-7.34617e-11               lu0_ss=2.87957e-11                lu0_mc=1.20418e-10 wu0_ff=5.26829e-11                wu0_ss=-2.10731e-10               wu0_mc=8.42924e-10 pu0_ff=-4.10925e-18               pu0_ss=1.6437e-17                 pu0_mc=-6.57481e-17 vsat_ff=-11108.8                   vsat_fs=-3817.59                   vsat_ss=5445.31 vsat_mc=-5789.31                   lvsat_ff=0.000866484                lvsat_fs=0.000297772 lvsat_ss=-0.000424734               lvsat_mc=0.000451566                wvsat_ff=0.00400389 wvsat_fs=0.00105365                 wvsat_ss=-0.00400389                wvsat_mc=0.00316096 pvsat_ff=-3.12303e-10               pvsat_fs=-8.21851e-11               pvsat_ss=3.12303e-10 pvsat_mc=-2.46555e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.16 nmos ( level=54                         lmin=9e-007                     lmax=9.019e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.45754533 lvth0=1.1681876e-008             wvth0=2.2421495e-009             pvth0=-4.7762897e-016 k2=-0.027815835               lk2=-4.8707545e-009            wk2=-1.3990834e-009 pk2=8.1662687e-017             cit=0.0012661442               lcit=2.762697e-010 wcit=1.0725706e-010             pcit=-1.1807325e-016            voff=-0.21173496 lvoff=-1.0122674e-008            wvoff=5.9214613e-009             pvoff=-1.3488448e-016 eta0=0.0065925926               weta0=3.8844444e-010             etab=-0.032464815 wetab=-1.7140111e-009            u0=0.023288578                lu0=9.3954323e-010 wu0=-1.2696989e-010            pu0=1.4617382e-016             ua=-1.1726588e-009 lua=7.0017383e-017             wua=-2.8632273e-018            pua=-1.8213062e-023 ub=1.7561513e-018             lub=-1.6261115e-025            wub=-2.8970265e-027 pub=2.6387608e-032             uc=1.0162419e-010             luc=-2.4807598e-017 wuc=-2.2683707e-018            puc=3.0741358e-024             vsat=86148.148 a0=1.0477386                  la0=5.3427713e-007             wa0=8.1808091e-008 pa0=2.5960026e-014             ags=0.4758665                  lags=6.8069412e-007 wags=2.5360847e-008             pags=-1.6092928e-014            keta=-0.0010528601 lketa=-4.5630004e-008            wketa=-1.2158006e-009            pketa=1.3264346e-015 pclm=1.1857887                  lpclm=1.277307e-007              wpclm=-2.129251e-009 ppclm=1.9137708e-014             pdiblc2=0.00065510221              lpdiblc2=5.3885136e-009 wpdiblc2=-5.4891665e-011            ppdiblc2=2.6605498e-016             agidl=1.5653042e-010 lagidl=-5.7917244e-018            wagidl=-5.6236941e-018            pagidl=2.8486722e-024 aigbacc=0.013531                   aigc=0.01140553                 laigc=-4.478835e-011 waigc=-4.8961103e-012            paigc=2.3646935e-018             aigsd=0.010858092 laigsd=-6.9758596e-011            waigsd=-1.8007144e-012            paigsd=9.3021702e-018 tvoff=0.00153441                 ltvoff=-1.95787e-010              wtvoff=6.91307e-011 ptvoff=2.63602e-017               kt1=-0.13314488                lkt1=-2.6296896e-008 wkt1=-3.6460274e-009            pkt1=2.7433063e-015             kt2=-0.065031111 lkt2=3.9414044e-009             ute=-0.54343799                lute=-7.1522623e-008 wute=-3.007877e-008             pute=1.4205921e-014             ua1=1.7025024e-009 lua1=-1.3557722e-016            wua1=6.7979794e-018             pua1=-1.1116387e-024 ub1=-4.8698738e-019            lub1=-9.4627282e-026            wub1=-8.6409892e-026 pub1=2.3256143e-032             uc1=3.8578041e-010             luc1=-6.3938339e-017 wuc1=-1.449502e-017             puc1=4.59305e-024               at=121939.87 lat=-0.017435527               wat=-0.00022114486             pat=1.98765e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-3.8844444e-010            pkt2=3.8120744e-030             lvsat=0 wvsat=0.0027191111               pvsat=0                          vth0_mcl=-7.69662e-05 lvth0_mcl=6.93235e-10                wvth0_mcl=2.12427e-11                pvth0_mcl=-1.91333e-16 cit_mcl=7.69662e-06                lcit_mcl=-6.93235e-11               wcit_mcl=-2.12427e-12 pcit_mcl=1.91333e-17                ags_ff=0.113403                   ags_ss=-0.170104 ags_sf=-0.113403                  lags_ff=-1.00701e-07               lags_ss=1.51052e-07 lags_sf=1.00701e-07                wags_ff=-1.29279e-08               wags_ss=1.93918e-08 wags_sf=1.29279e-08                pags_ff=1.148e-14                  pags_ss=-1.722e-14 pags_sf=-1.148e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.17 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.46515984 lvth0=4.920192e-009              wvth0=1.9302706e-009             pvth0=-2.0068054e-016 k2=-0.036349348               lk2=2.7070047e-009             wk2=-5.4815355e-010 pk2=-6.7396298e-016            cit=0.0010004118               lcit=5.1224004e-010 wcit=8.3824615e-012             pcit=-3.0272612e-017            voff=-0.22213383 lvoff=-8.8847624e-010            wvoff=6.5256763e-009             pvoff=-6.7142739e-016 eta0=0.0065925926               weta0=3.8844444e-010             etab=-0.032464815 wetab=-1.7140111e-009            u0=0.024921132                lu0=-5.1016443e-010 wu0=-1.8111528e-011            pu0=4.9507594e-017             ua=-9.5892905e-010 lua=-1.1977467e-016            wua=-1.9463958e-017            pua=-3.4716135e-024 ub=1.590703e-018              lub=-1.5693068e-026            wub=2.7609477e-026 pub=-7.0216727e-034            uc=7.5132791e-011             luc=-1.283234e-018 wuc=4.3190767e-018             puc=-2.7755176e-024            vsat=86148.148 a0=1.160356                   la0=4.3427293e-007             wa0=2.721945e-007 pa0=-1.4310311e-013            ags=0.7326681                  lags=4.526543e-007 wags=5.1916755e-008             pags=-3.9674574e-014            keta=-0.03534432 lketa=-1.5179188e-008            wketa=5.4845248e-010             pketa=-2.4022219e-016 pclm=1.2322963                  lpclm=8.6432e-008                wpclm=1.9422222e-008 ppclm=-5.0058424e-029            pdiblc2=0.007326278                lpdiblc2=-5.3549053e-010 wpdiblc2=1.9909569e-010             ppdiblc2=4.051421e-017              agidl=1.6505449e-010 lagidl=-1.3361097e-017            wagidl=-3.8059943e-018            pagidl=1.2345547e-024 aigbacc=0.013531                   aigc=0.011391469                laigc=-3.2301514e-011 waigc=-4.2079855e-012            paigc=1.7536388e-018             aigsd=0.010752106 laigsd=2.4356448e-011             waigsd=2.1674299e-011             paigsd=-1.1543641e-017 tvoff=0.00118368                 ltvoff=1.1566e-010                wtvoff=1.29016e-010 ptvoff=-2.68183e-017              kt1=-0.17363761                lkt1=9.6606471e-009 wkt1=1.3021815e-009             pkt1=-1.6507033e-015            kt2=-0.074435556 lkt2=1.2292551e-008             ute=-0.60728954                lute=-1.4822448e-008 wute=-1.8688088e-008            pute=4.0909956e-015             ua1=2.1728384e-009 lua1=-5.5323566e-016            wua1=-5.4878196e-017            pua1=5.3656805e-023 ub1=-1.1943955e-018            lub1=5.3355114e-025             wub1=4.9803757e-027 pub1=-5.7898415e-032            uc1=3.417521e-010              luc1=-2.4841197e-017 wuc1=-6.2979793e-018            puc1=-2.6859224e-024            at=163801.69 lat=-0.054608825               wat=0.0017848236               pat=2.0635005e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=7.4581333e-010             pkt2=-1.0072209e-015            lvsat=0 wvsat=0.0027191111               pvsat=0                          vth0_mcl=0.000703702 lvth0_mcl=1.9e-16                    wvth0_mcl=-1.94222e-10               pvth0_mcl=-1.5e-22 cit_mcl=-0.000138864               lcit_mcl=6.08225e-11                wcit_mcl=3.83265e-11 pcit_mcl=-1.6787e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.18 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.48188123 lvth0=-2.4037755e-009            wvth0=-2.3545728e-010            pvth0=7.4790828e-016 k2=-0.028878356               lk2=-5.6528987e-010            wk2=-3.248966e-009 pk2=5.0899286e-016             cit=0.0021631207               lcit=2.9735547e-012 wcit=-1.1416869e-010            pcit=2.3404792e-017             voff=-0.21494454 lvoff=-4.0373858e-009            wvoff=5.185462e-009              pvoff=-8.4413523e-017 eta0=0.0065925926               weta0=3.8844444e-010             etab=-0.032464815 wetab=-1.7140111e-009            u0=0.025829923                lu0=-9.0821491e-010 wu0=1.085865e-010              pu0=-5.9861414e-018            ua=-1.0945937e-009 lua=-6.0353564e-017            wua=-1.7325991e-017            pua=-4.4080431e-024 ub=1.7010773e-018             lub=-6.4037014e-026            wub=1.4864972e-026 pub=4.879926e-033              uc=1.2269436e-010             luc=-2.21152e-017 wuc=-7.29288e-018              puc=2.3105195e-024             vsat=83205.989 a0=3.2399527                  la0=-4.7659043e-007            wa0=-5.2956176e-008 pa0=-6.8711137e-016            ags=1.6671241                  lags=4.3362559e-008 wags=1.8986271e-008             pags=-2.5251022e-014            keta=-0.016980988 lketa=-2.3222327e-008            wketa=-2.6024782e-009            pketa=1.1398854e-015 pclm=1.4780627                  lpclm=-2.1213675e-008            wpclm=-5.9760684e-009 ppclm=1.1124451e-014             pdiblc2=0.0023769213               lpdiblc2=1.6323277e-009 wpdiblc2=3.8038754e-010             ppdiblc2=-3.8891618e-017            agidl=1.3810376e-010 lagidl=-1.5566803e-018            wagidl=-1.5724321e-018            pagidl=2.5625448e-025 aigbacc=0.013531                   aigc=0.011328174                laigc=-4.578474e-012 waigc=3.7670496e-012             paigc=-1.7394266e-018            aigsd=0.010831893 laigsd=-1.0589997e-011            waigsd=-1.039402e-011             paigsd=2.5022822e-018 tvoff=0.00184278                 ltvoff=-1.73027e-010              wtvoff=4.41201e-011 ptvoff=1.03662e-017               kt1=-0.11908538                lkt1=-1.4233228e-008 wkt1=-4.1959721e-009            pkt1=7.5748799e-016             kt2=-0.04637037 ute=-0.51341182                lute=-5.5940886e-008            wute=-2.8691254e-008 pute=8.4723821e-015             ua1=9.5169365e-010             lua1=-1.8374239e-017 wua1=1.0532586e-016             pua1=-1.6512572e-023            ub1=5.6208724e-019 lub1=-2.357883e-025             wub1=-2.2447308e-025            pub1=4.2602199e-032 uc1=4.4854701e-010             luc1=-7.1617368e-017            wuc1=-2.8685128e-017 puc1=7.1196488e-024             at=30761.504                  lat=0.0036627767 wat=0.0045634803               pat=-1.0107016e-009 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-1.5537778e-009            lvsat=0.0012886659               wvsat=0.0031153637 pvsat=-1.7355865e-010            vth0_mcl=-0.000168091               lvth0_mcl=3.81846e-10 wvth0_mcl=-1.94222e-10               pvth0_mcl=9e-24                      vsat_ff=742.64 lvsat_ff=-0.000325276               wvsat_ff=-8.4661e-05                pvsat_ff=3.70815e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.19 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.46588846 lvth0=8.5874893e-010             wvth0=3.7521165e-009             pvth0=-6.5556762e-017 k2=-0.03875208                lk2=1.4489498e-009             wk2=-1.3083903e-009 pk2=1.1311543e-016             cit=0.00077207585              lcit=2.867467e-010 wcit=3.3135822e-012             pcit=-5.6159151e-019            voff=-0.22004808 lvoff=-2.9962628e-009            wvoff=5.4594716e-009             pvoff=-1.4031148e-016 eta0=0.0065925926               weta0=3.8844444e-010             etab=-0.032464815 wetab=-1.7140111e-009            u0=0.018135386                lu0=6.6147054e-010 wu0=6.4698197e-010             pu0=-1.1581882e-016            ua=-1.6689509e-09 lua=5.6815303e-17              wua=-1.743237e-17              pua=-4.3863419e-24 ub=1.6309009e-018             lub=-4.9721024e-026            wub=3.7535757e-026 pub=2.5508592e-034             uc=1.6710794e-011             luc=-4.94553e-019 wuc=5.5680737e-018             puc=-3.1311508e-025            vsat=76710.998 a0=2.6229134                  la0=-3.5071441e-007            wa0=-1.9386881e-007 pa0=2.8059067e-014             ags=1.8052054                  lags=1.5193979e-008 wags=-1.6966526e-007            pags=1.323389e-014              keta=-0.087299859 lketa=-8.8772777e-009            wketa=1.2261896e-009             pketa=3.5883721e-016 pclm=1.2172487                  lpclm=3.1992381e-008             wpclm=9.1839365e-008 ppclm=-8.8298971e-015            pdiblc2=0.018231683                lpdiblc2=-1.6020437e-009 wpdiblc2=-3.8388765e-010            ppdiblc2=1.1702052e-016             agidl=1.3846782e-010 lagidl=-1.6309476e-018            wagidl=-4.2949959e-019            pagidl=2.3096239e-026 aigbacc=0.013531                   aigc=0.011359905                laigc=-1.1051623e-011 waigc=-5.2371403e-012            paigc=9.7428104e-020             aigsd=0.010808616 laigsd=-5.8415529e-012            waigsd=1.0873671e-011             paigsd=-1.8363267e-018 tvoff=0.000610087                ltvoff=7.84431e-011               wtvoff=1.64278e-010 ptvoff=-1.41461e-017              kt1=-0.20549148                lkt1=3.3936163e-009 wkt1=2.6711891e-009             pkt1=-6.434129e-016             kt2=-0.041784833 lkt2=-9.3544973e-010            ute=-0.85735633                lute=1.4223794e-008 wute=2.0788622e-008             pute=-1.6215125e-015            ua1=1.23071e-009 lua1=-7.5293573e-017            wua1=6.7742203e-017             pua1=-8.8455058e-024 ub1=-1.0618004e-018            lub1=9.5484769e-026             wub1=-5.3227155e-026 pub1=7.6680298e-033             uc1=2.3654321e-011             luc1=1.5060741e-017 wuc1=1.4631407e-017             puc1=-1.7169244e-024            at=49028.188 lat=-6.3626953e-005            wat=-0.0021256581              pat=3.5388265e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-1.7942434e-009            pkt2=4.9054984e-017             lvsat=0.0026136441 wvsat=0.0013610886               pvsat=1.8431348e-010             vth0_mcl=0.00170371 lvth0_mcl=4.4e-16                    wvth0_mcl=-1.94222e-10               pvth0_mcl=8e-24 vsat_ff=-1379.19                   lvsat_ff=0.000107577                wvsat_ff=0.000157228 pvsat_ff=-1.22637e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_12_mac.20 nmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.44023233 lvth0=2.859927e-009              wvth0=1.5397561e-009             pvth0=1.0700735e-016 k2=-0.041021734               lk2=1.6259828e-009             wk2=-2.4527158e-010 pk2=3.0192166e-017             cit=0.00076465916              lcit=2.8732521e-010 wcit=2.8991369e-010             pcit=-2.29164e-017              voff=-0.22126407 lvoff=-2.9014158e-009            wvoff=6.0357917e-009             pvoff=-1.8526445e-016 eta0=0.0065925926               weta0=3.8844444e-010             etab=-0.032465093 wetab=-1.7139794e-009            u0=0.022902432                lu0=2.8964096e-010 wu0=-4.2295126e-010            pu0=-3.2364026e-017            ua=-1.3845631e-09 lua=3.4633054e-17              wua=-1.1314933e-16             pua=3.0795806e-24 ub=1.1276014e-018             lub=-1.0463668e-026            wub=1.2813444e-025 pub=-6.8116116e-033            uc=5.0534979e-012             luc=4.1471605e-019 wuc=3.0212346e-018             puc=-1.1446163e-025            vsat=50592.672 a0=-8.00553                   la0=4.7830417e-007             wa0=1.4556078e-006 pa0=-1.0060011e-013            ags=-1.9409358                 lags=3.0739299e-007 wags=3.7915415e-007             pags=-2.9574024e-014            keta=-0.52292181 lketa=2.5101235e-008             wketa=4.2513086e-008             pketa=-2.8615407e-015 pclm=1.0915226                  lpclm=4.1799012e-008             wpclm=4.8339753e-008 ppclm=-5.4369274e-015            pdiblc2=-0.010870335               lpdiblc2=6.6791372e-010 wpdiblc2=2.0726264e-009             ppdiblc2=-7.4587575e-017            agidl=1.2209221e-010 lagidl=-3.5364999e-019            wagidl=-6.9460837e-018            pagidl=5.313898e-025 aigbacc=0.026768361                aigc=0.011427229                laigc=-1.6302862e-011 waigc=-5.1480866e-012            paigc=9.0481918e-020             aigsd=0.010590078 laigsd=1.1204423e-011             waigsd=-1.3516032e-011            paigsd=6.6070114e-020 tvoff=0.000680132                ltvoff=7.29796e-011               wtvoff=9.08988e-011 ptvoff=-8.42245e-018              kt1=-0.18703356                lkt1=1.953898e-009 wkt1=-1.7012958e-008            pkt1=8.9195055e-016             kt2=-0.054544737 lkt2=5.982279e-011              ute=-0.8130316                 lute=1.0766465e-008 wute=-5.491957e-009             pute=4.2837265e-016             ua1=4.727019e-010 lua1=-1.6168942e-017            wua1=1.4844662e-017             pua1=-4.7194975e-024 ub1=2.2589226e-019             lub1=-4.9552565e-027            wub1=-5.3374425e-026 pub1=7.6795169e-033             uc1=1.4090535e-010             luc1=5.9151605e-018 wuc1=-1.2516543e-017            puc1=4.006157e-025              at=28114.31 lat=0.0015676555               wat=0.0073190406               pat=-3.8280385e-010 jtsswgs='2e-007*(1+21*0.3*iboffn_flag_12)'                                 jtsswgd='2e-007*(1+21*0.3*iboffn_flag_12)' wkt2=-9.5365269e-010            pkt2=-1.651109e-017             lvsat=0.0046508734 wvsat=0.0086131138               pvsat=-3.8134449e-010            letab=2.1662365e-014 petab=-2.4695097e-021            laigbacc=-1.0325142e-009            waigbacc=-1.5090592e-009 paigbacc=1.1770662e-016             vth0_mcl=-0.0100427                 lvth0_mcl=9.16222e-10 wvth0_mcl=2.00572e-09                pvth0_mcl=-1.71595e-16               cit_mcl=-0.000489431 lcit_mcl=3.81758e-11                wcit_mcl=-7.33309e-11               pcit_mcl=5.71982e-18 voff_mcl=0.00377564                 lvoff_mcl=-2.94499e-10               wvoff_mcl=-7e-17 pvoff_mcl=-8e-24                     u0_ss=-0.00192977                u0_ff=0.00192977 u0_mc=0.00124456                 lu0_ss=1.50522e-10                lu0_ff=-1.50522e-10 lu0_mc=-9.70757e-11               wu0_ss=2.19994e-10                wu0_ff=-2.19994e-10 wu0_mc=7.33315e-11                pu0_ss=-1.71595e-17               pu0_ff=1.71595e-17 pu0_mc=-5.7198e-18                vsat_ss=-15438.2                   vsat_ff=5789.31 vsat_mc=9648.85                    lvsat_ss=0.00120418                 lvsat_ff=-0.000451566 lvsat_mc=-0.000752611               wvsat_ss=0.00175995                 wvsat_ff=-0.000659982 wvsat_mc=-0.00109997                pvsat_ss=-1.37276e-10               pvsat_ff=5.14786e-11 pvsat_mc=8.57976e-11 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model pch_12_mac.global pmos ( modelid=8                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_12'              permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=2.687e-009                 toxm=2.687e-009                 dtox=4.2747e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=-1.2e-008 xw=6e-009                     dlc=8e-009                     dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.47263 k3=-1.7282                    k3b=1.7496                     w0=0 dvt0=2.5                        dvt1=0.62                       dvt2=0 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.47671                    minv=-0.38                      voffl=0 dvtp0=4.5308e-007                dvtp1=0.1                        lpe0=5e-009 lpeb=6e-009                     xj=8.5e-008                   ngate=1.47e+020 ndep=6e+017                     nsd=1e+020                     phin=0.2 cdsc=0                          ud=0                          cdscb=0 cdscd=0                          nfactor=0.7                        a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=0.3 delta=0.014                      pscbe1=9.264e+008                 pscbe2=1e-020 fprout=0                          pdits=0                          pditsd=0 pditsl=0                          rsh=16.7                       rdsw=100.05 prwg=0                          prwb=0                          wr=1 alpha0=1.8425e-006                alpha1=8                          beta0=19 bgidl=1e+009                     cgidl=6.3146                     egidl=0.020298 aigbacc=0.011638                   bigbacc=0.0042384                  cigbacc=0.245 nigbacc=3.3599                     aigbinv=0.012555658                bigbinv=0.0032277133 cigbinv=0.006                      eigbinv=1.1                        nigbinv=3.0379743 bigc=0.0015262                  cigc=0.21515                    bigsd=0.00033025956 cigsd=0.0011                     nigc=1.9562914                  poxedge=1 pigcd=3.3707624                  ntox=1                          vfbsdoff=0.01 cgso=9.2e-011                   cgdo=9.2e-011                   cgbo=0 cgdl=1e-011                     cgsl=1e-011                     clc=0 cle=0.6                        cf='9.1e-011+8.7e-11*ccoflag_12' ckappas=0.6                        ckappad=0.6                        acde=0.37295 moin=5                          noff=2.4263                     voffcv=-0.133 tvfbsdoff=0.1                        kt1l=0                          prt=0 fnoimod=1.000000e+00               tnoimod=0                          em=1.000000e+07 ef=1.200000e+00               noia=0                          noib=0 noic=0                          jss=4.90e-07                   jsd=4.90e-07 jsws=1.01e-13                   jswd=1.01e-13                   jswgs=1.01e-13 jswgd=1.01e-13                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=7.42                       bvd=7.42 xjbvs=1                          xjbvd=1                          njtsswg=11 xtsswgs=0.55                       xtsswgd=0.55                       tnjtsswg=2 vtsswgs=8                          vtsswgd=8                          pbs=0.816 pbd=0.816                      cjs=0.001878                   cjd=0.001878 mjs=0.449                      mjd=0.449                      pbsws=0.742 pbswd=0.742                      cjsws=1.13e-010                  cjswd=1.13e-010 mjsws=0.253                      mjswd=0.253                      pbswgs=0.91 pbswgd=0.91                       cjswgs=1.86e-010                  cjswgd=1.86e-010 mjswgs=0.71                       mjswgd=0.71                       tpb=0.00100 tcj=0.00075                    tpbsw=0.00098                    tcjsw=0.00041 tpbswg=0.00125                    tcjswg=0.0010                     xtis=3 xtid=3                          dmcg=4.2e-008                   dmci=4.2e-008 dmdg=0                          dmcgt=0                          dwj=0 xgw=0                          xgl=-5.1e-009                  rshg=14.4 gbmin=1e-012                     rbpb=50                         rbpd=50 rbps=50                         rbdb=50                         rbsb=50 ngcon=1                          xrcrg1=12                         xrcrg2=1 k2we=0                          ku0we=-0.00055                   kvth0we=-0.0008 lk2we=0                          lku0we=-4.5e-11                   lkvth0we=2.5e-011 pk2we=0                          pku0we=1.8e-17                    pkvth0we=-2.178e-018 scref=1e-6                       web=1467.2                     wec=-6232.7 wk2we=0                          wku0we=-3e-10                     wkvth0we=4e-011 wpemod=1                          lintnoi=-1.5e-08 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.11 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.6 iboffn_flag='iboffn_flag_12' iboffp_flag='iboffp_flag_12' sigma_factor='sigma_factor_12' ccoflag='ccoflag_12' rcoflag='rcoflag_12' rgflag='rgflag_12' mismatchflag='mismatchflag_mos_12' globalflag='globalflag_mos_12' totalflag='totalflag_mos_12' global_factor='global_factor_12' local_factor='local_factor_12' sigma_factor_flicker='sigma_factor_flicker_12' noiseflag='noiseflagp_12' noiseflag_mc='noiseflagp_12_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w11='2.3875*0.35355' w12='0.70711*0.35355' w13='0.54772*0.32451' w14='0.54772*-0.16328' w15='0.54772*0.12195' w16='0.54772*0.66871' w17='0.54772*0.32929' w18='0.54772*-0.21807' w19='0' w20='0' tox_c='toxp_12'                  dxl_c='dxlp_12'                  dxw_c='dxwp_12' cj_c='cjp_12'                   cjsw_c='cjswp_12'                 cjswg_c='cjswgp_12' cgo_c='cgop_12'                  cgl_c='cglp_12'                  ddlc_c='ddlcp_12' ntox_c='ntoxp_12'                 cf_c='cfp_12'                   dvth_c='dvthp_12' dlvth_c='dlvthp_12'                dwvth_c='dwvthp_12'                dpvth_c='dpvthp_12' du0_c='du0p_12'                  dlu0_c='dlu0p_12'                 dwu0_c='dwu0p_12' dpu0_c='dpu0p_12'                 dvsat_c='dvsatp_12'                dlvsat_c='dlvsatp_12' dwvsat_c='dwvsatp_12'               dpvsat_c='dpvsatp_12'               dk2_c='dk2p_12' dlk2_c='dlk2p_12'                 dwk2_c='dwk2p_12'                 dpk2_c='dpk2p_12' dvoff_c='dvoffp_12'                dlvoff_c='dlvoffp_12'               dwvoff_c='dwvoffp_12' dpvoff_c='dpvoffp_12'               dags_c='dagsp_12'                 dlags_c='dlagsp_12' dwags_c='dwagsp_12'                dpags_c='dpagsp_12'                dcit_c='dcitp_12' dlcit_c='dlcitp_12'                dwcit_c='dwcitp_12'                dpcit_c='dpcitp_12' deta0_c='deta0p_12'                dpclm_c='dpclmp_12'                dua1_c='dua1p_12' dlua1_c='dlua1p_12'                dwua1_c='dwua1p_12'                dpua1_c='dpua1p_12' duc_c='ducp_12'                  dluc_c='dlucp_12'                 dwuc_c='dwucp_12' dpuc_c='dpucp_12'                 dketa_c='dketap_12'                dlketa_c='dlketap_12' dwketa_c='dwketap_12'               dpketa_c='dpketap_12'               jtsswg_c='jtsswgp_12' ss_flag_c='ss_flagp_12'              ff_flag_c='ff_flagp_12'              sf_flag_c='sf_flagp_12' fs_flag_c='fs_flagp_12'              monte_flag_c='monte_flagp_12'          c1f_c='c1fp_12' c2f_c='c2fp_12'                  c3f_c='c3fp_12' global_mc='global_mc_flag_12' tox_g='toxp_12_ms_global'        dxl_g='dxlp_12_ms_global'        dxw_g='dxwp_12_ms_global' cj_g='cjp_12_ms_global'         cjsw_g='cjswp_12_ms_global'       cjswg_g='cjswgp_12_ms_global' cgo_g='cgop_12_ms_global'        cgl_g='cglp_12_ms_global'        ntox_g='ntoxp_12_ms_global' cf_g='cfp_12_ms_global'         dvth_g='dvthp_12_ms_global'       dlvth_g='dlvthp_12_ms_global' dwvth_g='dwvthp_12_ms_global'      dpvth_g='dpvthp_12_ms_global'      du0_g='du0p_12_ms_global' dlu0_g='dlu0p_12_ms_global'       dwu0_g='dwu0p_12_ms_global'       dpu0_g='dpu0p_12_ms_global' dvsat_g='dvsatp_12_ms_global'      dwvsat_g='dwvsatp_12_ms_global' dpvsat_g='dpvsatp_12_ms_global'     dk2_g='dk2p_12_ms_global'        dlk2_g='dlk2p_12_ms_global' dwk2_g='dwk2p_12_ms_global'       dpk2_g='dpk2p_12_ms_global'       dlvoff_g='dlvoffp_12_ms_global' dpvoff_g='dpvoffp_12_ms_global'     dags_g='dagsp_12_ms_global'       dwags_g='dwagsp_12_ms_global' dcit_g='dcitp_12_ms_global'       dlcit_g='dlcitp_12_ms_global'      dwcit_g='dwcitp_12_ms_global' dpcit_g='dpcitp_12_ms_global'      deta0_g='deta0p_12_ms_global'      dpclm_g='dpclmp_12_ms_global' dua1_g='dua1p_12_ms_global'       dluc_g='dlucp_12_ms_global'       dlketa_g='dlketap_12_ms_global' ss_flag_g='ss_flagp_12_ms_global'    ff_flag_g='ff_flagp_12_ms_global' monte_flag_g='monte_flagp_12_ms_global'                                        sf_flag_g='sf_flagp_12_ms_global' fs_flag_g='fs_flagp_12_ms_global' weight1=-3.4730769 weight2=2.2129371 weight3=1.5223776 weight4=-0.6993007 weight5=-0.48693706 tox_1=4.3342957e-012 tox_2=-9.6864903e-012 tox_3=-2.1640978e-013 tox_4=3.7476963e-011 tox_5=7.5517924e-013 dxl_1=2.1262979e-010 dxl_2=-4.7518952e-010 dxl_3=-1.0616989e-011 dxl_4=-1.8384982e-009 dxl_5=3.7046963e-011 dxw_1=-7.1356929e-010 dxw_2=-8.0891919e-010 dxw_3=-9.5014905e-012 dxw_4=5.993894e-025 dxw_5=-5.9015941e-009 cj_1=1.3034e-005 cj_2=-3.5938e-006 cj_3=-1.7529e-007 cj_4=6.1114e-021 cj_5=-1.0826e-006 cjsw_1=7.8426e-013 cjsw_2=-2.1624e-013 cjsw_3=-1.0547e-014 cjsw_4=-7.2349e-028 cjsw_5=-6.5141e-014 cjswg_1=1.2909e-012 cjswg_2=-3.5594e-013 cjswg_3=-1.7361e-014 cjswg_4=-1.0066e-028 cjswg_5=-1.0722e-013 cgo_1=-6.3851e-013 cgo_2=1.7606e-013 cgo_3=8.587e-015 cgo_4=1.0263e-027 cgo_5=5.3035e-014 cgl_1=-6.9404e-014 cgl_2=1.9137e-014 cgl_3=9.3337e-016 cgl_4=-3.2542e-029 cgl_5=5.7647e-015 ntox_1=-0.31727 ntox_2=0.087481 ntox_3=0.0042668 ntox_4=-1.4519e-016 ntox_5=0.026353 cf_1=-6.3157e-013 cf_2=1.7414e-013 cf_3=8.4937e-015 cf_4=-2.8903e-028 cf_5=5.2459e-014 dvth_1=-0.0032683 dvth_2=-0.0039068 dvth_3=0.00013258 dvth_4=-1.5551e-018 dvth_5=0.00090272 dlvth_1=-1.1841e-010 dlvth_2=-1.1154e-010 dlvth_3=-1.9536e-012 dlvth_4=3.08e-026 dlvth_5=2.8772e-011 dwvth_1=-1.248e-010 dwvth_2=2.4577e-012 dwvth_3=2.0274e-011 dwvth_4=-1.8533e-025 dwvth_5=1.3521e-011 dpvth_1=-3.1918e-017 dpvth_2=-1.5174e-017 dpvth_3=-8.5744e-019 dpvth_4=-2.5116e-032 dpvth_5=5.5964e-018 du0_1=5.8079e-005 du0_2=0.00012922 du0_3=6.2603e-006 du0_4=-4.3061e-020 du0_5=-2.5026e-005 dlu0_1=-3.5371e-013 dlu0_2=2.736e-011 dlu0_3=-2.4653e-012 dlu0_4=6.4673e-028 dlu0_5=-3.5478e-012 dwu0_1=1.095e-012 dwu0_2=2.231e-011 dwu0_3=-2.7648e-012 dwu0_4=-2.8754e-027 dwu0_5=-3.0031e-012 dpu0_1=4.8652e-019 dpu0_2=2.298e-018 dpu0_3=1.9417e-019 dpu0_4=1.5154e-034 dpu0_5=-4.8256e-019 dvsat_1=665.76 dvsat_2=742.19 dvsat_3=115.01 dvsat_4=-5.3235e-013 dvsat_5=-189.57 dwvsat_1=0.00010571 dwvsat_2=0.00013055 dwvsat_3=6.2323e-005 dwvsat_4=-7.7939e-020 dwvsat_5=-2.9819e-005 dpvsat_1=8.6842e-013 dpvsat_2=7.7713e-012 dpvsat_3=1.375e-013 dpvsat_4=-2.3301e-027 dpvsat_5=-1.1242e-012 dk2_1=0.0015123 dk2_2=0.0011843 dk2_3=0.00011076 dk2_4=6.7634e-019 dk2_5=-0.00033603 dlk2_1=-7.7891e-012 dlk2_2=1.8211e-011 dlk2_3=-4.4578e-012 dlk2_4=3.3524e-027 dlk2_5=-1.4574e-012 dwk2_1=2.4771e-011 dwk2_2=-6.744e-012 dwk2_3=-1.046e-011 dwk2_4=1.0355e-026 dwk2_5=-2.0579e-012 dpk2_1=-5.6755e-018 dpk2_2=1.561e-018 dpk2_3=5.3204e-019 dpk2_4=8.7665e-034 dpk2_5=4.7143e-019 dlvoff_1=-1.492e-011 dlvoff_2=4.3721e-012 dlvoff_3=-3.018e-011 dlvoff_4=8.0247e-027 dlvoff_5=1.2381e-012 dpvoff_1=-1.2434e-018 dpvoff_2=3.6434e-019 dpvoff_3=-2.515e-018 dpvoff_4=4.7875e-034 dpvoff_5=1.0317e-019 dags_1=0.02711 dags_2=0.020875 dags_3=-0.0022904 dags_4=9.9746e-018 dags_5=-0.0063073 dwags_1=1.2171e-009 dwags_2=-3.3755e-009 dwags_3=-1.2235e-010 dwags_4=-1.339e-024 dwags_5=3.0228e-010 dcit_1=4.561e-006 dcit_2=-1.254e-006 dcit_3=-4.8302e-007 dcit_4=-1.845e-021 dcit_5=-3.7886e-007 dlcit_1=-1.983e-012 dlcit_2=5.4676e-013 dlcit_3=2.6668e-014 dlcit_4=-1.163e-027 dlcit_5=1.6471e-013 dwcit_1=-2.5012e-014 dwcit_2=1.6191e-014 dwcit_3=-1.0936e-012 dwcit_4=3.0228e-028 dwcit_5=2.0332e-015 dpcit_1=2.3599e-020 dpcit_2=-1.4761e-020 dpcit_3=9.7119e-019 dpcit_4=1.4464e-035 dpcit_5=-1.9207e-021 deta0_1=-0.0014872 deta0_2=0.00041007 deta0_3=2.0001e-005 deta0_4=-4.4644e-018 deta0_5=0.00012353 dpclm_1=-0.014872 dpclm_2=0.0041007 dpclm_3=0.00020001 dpclm_4=1.4097e-018 dpclm_5=0.0012353 dua1_1=7.9319e-012 dua1_2=-2.187e-012 dua1_3=-1.0667e-013 dua1_4=-3.8398e-027 dua1_5=-6.5882e-013 dluc_1=1.9766e-019 dluc_2=-5.1057e-020 dluc_3=-4.0773e-019 dluc_4=-2.8892e-034 dluc_5=-1.6434e-020 dlketa_1=-1.2848e-010 dlketa_2=3.3187e-011 dlketa_3=2.6503e-010 dlketa_4=4.8787e-026 dlketa_5=1.0682e-011 ss_flag_1=0.049735 ss_flag_2=-0.014574 ss_flag_3=0.1006 ss_flag_4=-5.004e-017 ss_flag_5=-0.0041269 ff_flag_1=-0.049414 ff_flag_2=0.012764 ff_flag_3=0.10193 ff_flag_4=8.6285e-017 ff_flag_5=0.0041084 monte_flag_1=0.0817808 monte_flag_2=-0.182765 monte_flag_3=-0.00408346 monte_flag_4=-0.707115 monte_flag_5=0.0142488 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.87 b_4=0.004                      c_4=0.001                      d_4=-0.00085 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=-0.0018                    mis_a_2=-0.1                       mis_a_3=0.05 mis_b_1=0.0021                     mis_b_2=0.05                       mis_b_3=0.05 mis_c_1=0.2922                     mis_c_2=0.0000                     mis_c_3=0.0000 mis_d_1=0.0005                     mis_d_2=0                          mis_d_3=0.25 mis_e_1=0.0033                     mis_e_2=-0.08                      mis_e_3=-0.05 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-1.2e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=60                         co_rsd=16.7                       bidirectionflag=1 designflag=1 cf0=9.1e-011                   cco=8.7e-11 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=1                          l_rjtsswg=0                          ll_rjtsswg=2 w_rjtsswg=0e-03                      ww_rjtsswg=2                          p_rjtsswg=0 noimod=1                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6               sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=1                   lreflod=0.9e-6              llodref=2 lod_clamp=-1e-90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=0 kvth00=-0e-9               lkvth00=0e-8                wkvth00=0e-8 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0e-11 lodeta00=1 wlod00=0 ku000=-1.0e-8             lku000=0.9e-15                  wku000=0.7e-15		   pku000=0 llodku000=1                   wlodku000=1 kvth000=-1.0e-9             lkvth000=0.08e-15	            wkvth000=0.15e-15		   pkvth000=-5.5e-24 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0.9e-6 ku01=-16.0e-8                lku01=0                wku01=-0e-15 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0.3 kvth01=0e-9                lkvth01=0e-24               wkvth01=-0.0e-19 pkvth01=0                   llodvth1=1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.00               lku02=2e-7              wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0 kvth02=2.5e-3             lkvth02=0                   wkvth02=0 pkvth02=0                   llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0e-4 lodeta02=1 wlod02=0 ku002=-0.010                   lku002=4e-10             wku002=0e-9         		pku002=0 llodku002=1                   wlodku002=1 kvth002=-0.001                 lkvth002=-13e-11             wkvth002=0e-10         	pkvth002=-1e-18 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0.2                lku03=-3e-9           wku03=-1.0e-8 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0.3 kvth03=0.005                lkvth03=0                   wkvth03=0 pkvth03=-1e-17              llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0.000 lodeta03=1 wlod03=0 ku003=0.00                   lku003=-1.5e5                   wku003=-1e-9         		pku003=0e-2 llodku003=-1                   wlodku003=1 kvth003=7.2e-3                   lkvth003=-1.5e-10             wkvth003=-3e-10         	pkvth003=0e-17 llodvth03=1                   wlodvth03=1                   steta003=0.0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=1 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='-0.05*1'              wkvth0dpl='-1e-8*1.5'                   wdplkvth0=1 lkvth0dpl='-1.0e-8*0'              ldplkvth0=1.0                 pkvth0dpl='-4.5e-15' ku0dpl=0.6                wku0dpl='2e-7*0.4'                   wdplku0=1 lku0dpl='-1.0e-7*0.5'              ldplku0=1.0                 pku0dpl='0.7e-14' keta0dpl=-0.2                wketa0dpl=0                   wdplketa0=1 kvsatdpl='1-0.5'                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=-3             ku0dpl_b2=-3 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx='1.0e-6*0'              wkvth0dpx=0                   wdpxkvth0=1 lkvth0dpx=0                   ldpxkvth0=1                   pkvth0dpx=0 ku0dpx=0                   wku0dpx=0                   wdpxku0=1 lku0dpx=0                   ldpxku0=1                   pku0dpx=0 keta0dpx=0                   wketa0dpx=0                   wdpxketa0=1 kvsatdpx=0                   wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps='-0.05*1.7'               wkvth0dps=0                   wdpskvth0=1 lkvth0dps='1.0e-7*1'             ldpskvth0=1.0                 pkvth0dps=0 ku0dps=4.5               wku0dps='-1.0e-8*5.5'                   wdpsku0=1 lku0dps='1.1e-8*2'        ldpsku0=1.2                 pku0dps='-1.0e-18*1*0' keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps='0.9'                 wdps=0 kvth0dps_b1=0.002            kvth0dps_b2=-0.000            dpsbinflg=1 ku0dps_b1=0.1                 ku0dps_b2=0.2 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa='0.002*1'               wkvth0dpa='-2.0e-9*0'            wdpakvth0=1 lkvth0dpa='-0.00e-7'            ldpakvth0=1.0                pkvth0dpa='6.0e-17*1' ku0dpa='-0.035'               wku0dpa='2e-9*0'               wdpaku0=1 lku0dpa='-4e-9*0'               ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa='1.10*1*0'                wdpa=0 kvth0dpa_b1=0.008             kvth0dpa_b2=0.000            dpabinflg=1 ku0dpa_b1=-0.08             ku0dpa_b2=-0.07 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1='0.0'                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2='-0.01*0'               wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2='-1.0e-9*0'              ldp2kvth0=1                   pkvth0dp2='-1e-16*1' ku0dp2=0.1                wku0dp2='2.0e-8*0'             wdp2ku0=1 lku0dp2=-0.0e-8              ldp2ku0=1.0                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=1.0                wdp2=0 kvth0dp2l='-0.03'              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l='3.0e-9'             ldp2lkvth0=1                  pkvth0dp2l='0e-15' ku0dp2l=0.57               wku0dp2l='-6.0e-8*1'            wdp2lku0=1 lku0dp2l=8e-10               ldp2lku0=1.2                pku0dp2l=-1e-17 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l='0.5'                wdp2l=0 kvth0dp2l_b1='0.016'            kvth0dp2l_b2='-0.016'           dp2lbinflg=1 ku0dp2l_b1='-0.08'            ku0dp2l_b2='0.06' keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a='0.005*0'              wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a='1.0e-9*0'             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=-0.00              wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a='-9.0e-5*0'            ldp2aku0='0.5*2'                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=0.010           kvth0dp2a_b2=-0.000           dp2abinflg=1 ku0dp2a_b1=-0.04              ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx=-0.020              wkvth0enx=-1.0e-9             wenxkvth0=1.0 lkvth0enx=-3.0e-8             lenxkvth0=1.0                 pkvth0enx=-0.85e-16 ku0enx=-1.8                wku0enx=-0.5e-7           wenxku0=1.0 lku0enx=0.1e-8             lenxku0=1.2                 pku0enx='-0.5e-16' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0.0                 wka0enx=0                   wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx=0.5                 wenx=0                   ku0enx0=-0.20 eny0=0.08e-6 enyref=0.08e-6             enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0.006               wkvth0eny='1e-9'              wenykvth0=1 lkvth0eny='1.0e-7*0'          lenykvth0=1.0                 pkvth0eny='4.0e-17*0' ku0eny='6.3'               wku0eny='1.0e-8*1.3'        wenyku0=1 ku0eny0='-0.11*-0'          wku0eny0='-1.0e-7*2.0'       weny0ku0=1 lku0eny='2.8e-4'            lenyku0=0.7                 pku0eny='0.0e-15' keta0eny=0e-4                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny='0.40'              weny=0 kvth0eny1='-6e-4*0'          wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1='3.0e-18*0' ku0eny1='-0.5e-3'          wku0eny1='-1.0e-9'          weny1ku0=1 lku0eny1='-0.6e-8'          leny1ku0=1.0                pku0eny1='-5.0e-18' keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1='1.0e-8*0'         weny1ka0=1 lka0eny1='4.0e-9*0'         leny1ka0=1.0                pka0eny1='3.0e-15*0' kvsateny1=0.50               weny1=0 rx_mode=1 rxref=1.8126e-5              ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=0.013               wkvth0rx=0e-9          	     wrxkvth0=1 lkvth0rx=-7e-9               lrxkvth0=1                	 pkvth0rx=0e-16 ku0rx=1.1              	 wku0rx=0.1e-8           	 wrxku0=1 lku0rx=4.2e-7        	     lrxku0=1                   pku0rx=-6e-16 keta0rx=0                	 wketa0rx=0                   wrxketa0=1 kvsatrx=1.9                 wrx=0                   ku0rx0=0.10 ry_mode=1 ryref=1.8027e-5           ringymax=0.9027e-5           ringymin=0.117e-6 kvth0ry=-0.010           	 wkvth0ry=-8.5e-9           	 wrykvth0=1 lkvth0ry=-5e-9               lrykvth0=1                 	 pkvth0ry=0 ku0ry=-0.9	          	 wku0ry=0           		 wryku0=1 lku0ry=0        			 lryku0=1      	         pku0ry=0 keta0ry=0                	 wketa0ry=0                   wryketa0=1 kvsatry=0.15                wry=0 kvth0ry0=0                	 ku0ry0=-0.00 sfxref=9.0e-8            sfxmax=1.53e-6            minwodx=0.0e-6 sfxmin=9.0e-8 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=0.0 kvth0odx1a=-0.011            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.07              lku0odx1a=1.6e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.6 kvth0odx1b=0.0003            lkvth0odx1b=1.8e-11           lodx1bkvth0=1.00 wkvth0odx1b=-0.0e-11           wodx1bkvth0=1.0               pkvth0odx1b=-0.7e-18 ku0odx1b=0.00245           lku0odx1b=0.8e-6           lodx1bku0=0.5 wku0odx1b=-0.0e-6           wodx1bku0=1.0               pku0odx1b=-1.0e-14 sfyref=7.92e-7 sfymin=0.144e-6 sfymax=1.53e-6           minwody=0.054e-6              wody=5e-7 kvth0odya=0                 lkvth0odya=0.0e-4            lodyakvth0=1.0 wkvth0odya=0.0e-7            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=0                 lku0odya=0.0e-6            lodyaku0=1.0 wku0odya=-0.0e-8           wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=-0.0e-2           wketa0ody=0                 wodyketa0=1 kvsatody=0.4 lrefody=1.0e-7            lodyref=1 kvth0odyb=0.020             lkvth0odyb=2.5e-9            lodybkvth0=1.0 wkvth0odyb=3.1e-8              wodybkvth0=1.0               pkvth0odyb=18e-16 ku0odyb=-0.35              lku0odyb=0e-9             lodybku0=0.9 wku0odyb=-3.0e-7           wodybku0=1.0               pku0odyb=-0.8e-13 web_mac=-4086.3  wec_mac=-7474.8 kvsatwe=0.3e-3 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model pch_12_mac.1 pmos ( level=54                         lmin=9e-007                     lmax=9.023e-06 wmin=9e-007                     wmax=1.351e-06                  vth0=-0.52939156 lvth0=8.5730835e-009             wvth0=8.7072411e-009             pvth0=-7.1927663e-015 k2=0.024496744                lk2=-1.0252889e-008            wk2=-2.348566e-008 pk2=9.2850183e-015             cit=0.00099042071              lcit=5.5849479e-010 wcit=-1.4908201e-010            pcit=2.7524705e-016             voff=-0.12973743 lvoff=-7.1763474e-009            wvoff=-3.1939024e-009            pvoff=-1.9857256e-015 eta0=0.06679608                 weta0=3.0082752e-008             etab=-0.14741947 wetab=2.6509077e-008             u0=0.01335196                 lu0=3.4013007e-009 wu0=-1.9249693e-009            pu0=2.6900874e-017             ua=1.7049273e-009 lua=1.8424761e-016             wua=-9.93491e-016              pua=1.6991216e-022 ub=1.8572786e-019             lub=1.1062405e-025             wub=5.7595657e-025 pub=-4.8660291e-032            uc=-3.2407504e-011            luc=1.5366222e-017 wuc=-1.2153244e-016            puc=3.940978e-023              vsat=90251.277 lvsat=0.044914143                wvsat=0.033721989                pvsat=-6.0903578e-008 a0=1.4190159                  la0=-7.2543478e-008            wa0=1.987226e-007 pa0=-1.2914079e-013            ags=0.56089065                 lags=1.9873219e-007 wags=-5.8716374e-008            pags=-1.5310627e-014            keta=-0.047328807 lketa=6.3474521e-008             wketa=6.3250015e-008             pketa=-7.7731957e-014 pclm=0.27158038                 lpclm=-1.3762968e-007            wpclm=6.1810145e-007 ppclm=-1.4740818e-013            pdiblc2=0.00021415901              lpdiblc2=2.5691388e-009 wpdiblc2=1.6461371e-010             ppdiblc2=-1.479548e-015             agidl=1.7487224e-010 lagidl=5.3308002e-017             wagidl=-2.0551274e-017            pagidl=-3.9973673e-023 aigc=0.0067795977               laigc=-4.4457234e-011            waigc=-5.2068405e-012 paigc=1.4828084e-017             aigsd=0.0061188628               laigsd=-1.2662126e-010 waigsd=-4.3338319e-011            paigsd=1.1588436e-016             tvoff=0.00149667 ltvoff=4.31948e-010               wtvoff=2.05769e-010               ptvoff=-8.66565e-016 kt1=-0.19783767                lkt1=-1.120789e-008             wkt1=9.7079897e-009 pkt1=-5.8031291e-015            kt2=-0.061606477               lkt2=-2.1186818e-009 wkt2=1.5637037e-009             pkt2=8.3976635e-015             ute=-0.78552888 lute=-2.0705761e-007            wute=-1.5197267e-007            pute=1.8074697e-013 ua1=2.9607486e-009             lua1=5.0560951e-016             wua1=-7.5483148e-016 pua1=-3.1873497e-022            ub1=-3.0661272e-018            lub1=-1.416941e-024 wub1=4.7160204e-025             pub1=1.1911685e-030             uc1=3.6392048e-010 luc1=1.2508854e-016             wuc1=7.352067e-017              puc1=-2.4444369e-022 at=128903.7                   lat=0.0098535111 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' u0_ff=0.000199677                u0_ss=-0.000199677               u0_sf=0.000110932 u0_fs=-0.000110932               lu0_ff=-1.77313e-10               lu0_ss=1.77313e-10 lu0_sf=-9.85072e-11               lu0_fs=9.85072e-11                wu0_ff=-1.6e-16 wu0_ss=1.6e-16                    wu0_sf=3.5e-16                    wu0_fs=-3.5e-16 pu0_ff=-1.2e-22                   pu0_ss=1.2e-22                    pu0_sf=-7e-23 pu0_fs=7e-23 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_12_mac.2 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=1.351e-06                  vth0=-0.51315929 lvth0=-5.8411681e-009            wvth0=5.0199765e-010             pvth0=9.3489838e-017 k2=0.022105782                lk2=-8.1297145e-009            wk2=-1.6778055e-008 pk2=3.3286652e-015             cit=0.0015964208               lcit=2.0366688e-011 wcit=3.4874881e-010             pcit=-1.6682672e-016            voff=-0.1228293 lvoff=-1.3310767e-008            wvoff=-5.5701903e-009            pvoff=1.2441794e-016 eta0=0.06679608                 weta0=3.0082752e-008             etab=-0.14741947 wetab=2.6509077e-008             u0=0.011487897                lu0=5.0565885e-009 wu0=5.6467955e-011             pu0=-1.7326154e-015            ua=1.502764e-009 lua=3.6376855e-016             wua=-3.3747604e-016            pua=-4.1262912e-022 ub=4.0541632e-019             lub=-8.44593e-026              wub=3.0761197e-025 pub=1.8962972e-031             uc=2.8544441e-011             luc=-3.8759105e-017 wuc=-1.4161762e-016            puc=5.7245418e-023             vsat=178250.42 lvsat=-0.033229096               wvsat=-0.055987037               pvsat=1.8758037e-008 a0=2.1455267                  la0=-7.1768507e-007            wa0=-4.1215767e-007 pa0=4.1332089e-013             ags=1.702142                   lags=-8.1469896e-007 wags=-1.122728e-006             pags=9.2953165e-013             keta=0.025807369 lketa=-1.4704031e-009            wketa=-2.2397711e-008            pketa=-1.6767764e-015 pclm=-0.18611207                lpclm=2.6880121e-007             wpclm=7.3058397e-007 ppclm=-2.4729266e-013            pdiblc2=0.0024279467               lpdiblc2=6.0329536e-010 wpdiblc2=-1.9001357e-009            ppdiblc2=3.5394941e-016             agidl=3.2979129e-010 lagidl=-8.4260119e-017            wagidl=-1.2873073e-016            pagidl=5.6089681e-023 aigc=0.0067743813               laigc=-3.9825062e-011            waigc=-1.8473952e-011 paigc=2.660928e-017              aigsd=0.0058513397               laigsd=1.1093921e-010 waigsd=2.3278565e-010             paigsd=-1.2931372e-016            tvoff=0.00287317 ltvoff=-7.90376e-010              wtvoff=-1.56853e-009              ptvoff=7.09012e-016 kt1=-0.1773809                 lkt1=-2.9373504e-008            wkt1=-2.3912388e-008 pkt1=2.4051766e-014             kt2=-0.0679575                 lkt2=3.5210268e-009 wkt2=1.2322122e-008             pkt2=-1.1558121e-015            ute=-0.47425552 lute=-4.8346836e-007            wute=-4.2981758e-007            pute=4.2747325e-013 ua1=4.874637e-009              lua1=-1.1939234e-015            wua1=-2.370496e-015 pua1=1.1159751e-021             ub1=-4.3720851e-018            lub1=-2.5725036e-025 wub1=1.3188767e-024             pub1=4.3878861e-031             uc1=9.7234185e-010 luc1=-4.1518963e-016            wuc1=-6.694597e-016             puc1=4.1532288e-022 at=107195.1                   lat=0.029130755 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=0.087301718                pat=-7.7523925e-008            vsat_ff=7795.3 vsat_ss=-2911.4                    vsat_sf=4866.7                     vsat_fs=-7795.3 lvsat_ff=-0.00692227                lvsat_ss=0.00258526                 lvsat_sf=-0.00432157 lvsat_fs=0.00692227                 wvsat_ff=-0.00265329                wvsat_ss=-0.00265335 wvsat_sf=6e-09                      wvsat_fs=0.00265329                 pvsat_ff=2.35616e-09 pvsat_ss=2.3562e-09                 pvsat_sf=-3.5e-14                   pvsat_fs=-2.35616e-09 ags_ff=0.0482351                  ags_ss=-0.341098                  ags_sf=0.585727 ags_fs=-0.194667                  lags_ff=-4.28328e-08               lags_ss=3.02895e-07 lags_sf=-5.20125e-07               lags_fs=1.72864e-07                wags_ff=1.32667e-07 wags_ss=1.32667e-07                wags_sf=-5.30668e-07               wags_fs=-2.4e-13 pags_ff=-1.17808e-13               pags_ss=-1.17809e-13               pags_sf=4.71233e-13 pags_fs=4e-19                      at_ff=14643.2                    at_sf=8785.9 at_ss=-14643.2                   at_fs=-8785.9                    lat_ff=-0.0130031 lat_sf=-0.00780188                lat_ss=0.0130031                  lat_fs=0.00780188 wat_ff=-0.0132667                 wat_sf=-0.00796002                wat_ss=0.0132667 wat_fs=0.00796002                 pat_ff=1.17808e-08                pat_sf=7.0685e-09 pat_ss=-1.17808e-08               pat_fs=-7.0685e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_12_mac.3 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=1.351e-06                  vth0=-0.51795864 lvth0=-3.7390554e-009            wvth0=2.7909679e-009             pvth0=-9.0907914e-016 k2=0.012252707                lk2=-3.8140674e-009            wk2=-7.1528791e-009 pk2=-8.8716194e-016            cit=0.00049820836              lcit=5.0138375e-010 wcit=4.5607979e-010             pcit=-2.1383769e-016            voff=-0.13464631 lvoff=-8.134918e-009             wvoff=-7.3767748e-009            pvoff=9.1570196e-016 eta0=0.06679608                 weta0=3.0082752e-008             etab=-0.14741947 wetab=2.6509077e-008             u0=0.019883386                lu0=1.3793641e-009 wu0=-6.2600954e-009            pu0=1.0340394e-015             ua=3.7910727e-009 lua=-6.3851066e-016            wua=-1.9447371e-015            pua=2.9135121e-022 ub=-2.8693609e-019            lub=2.1879106e-025             wub=8.5626822e-025 pub=-5.0681718e-032            uc=-1.6809573e-010            luc=4.7369288e-017 wuc=-1.400041e-018             puc=-4.1698822e-024            vsat=133194.1 lvsat=-0.01349443                wvsat=-0.031612767               pvsat=8.0821067e-009 a0=1.5595213                  la0=-4.6101468e-007            wa0=9.1732691e-007 pa0=-1.6899336e-013            ags=-3.474836                  lags=1.4528174e-006 wags=1.7296732e-006             pags=-3.1982007e-013            keta=0.12703627 lketa=-4.5808664e-008            wketa=-6.9796238e-008            pketa=1.9083779e-014 pclm=0.28734427                 lpclm=6.1427336e-008             wpclm=2.4976732e-007 ppclm=-3.6694963e-014            pdiblc2=0.0036356239               lpdiblc2=7.4332718e-011 wpdiblc2=-2.0440599e-009            ppdiblc2=4.1698822e-016             agidl=1.624527e-010 lagidl=-1.0965815e-017            wagidl=-2.9375794e-017            pagidl=1.2572221e-023 aigc=0.006584867                laigc=4.3182215e-011             waigc=1.5680205e-010 paigc=-5.0161608e-017            aigsd=0.0061476708               laigsd=-1.8853802e-011 waigsd=-1.3508979e-010            paigsd=3.1815722e-017             tvoff=0.00120263 ltvoff=-5.86815e-011              wtvoff=-2.3039e-010               ptvoff=1.22907e-016 kt1=-0.24517628                lkt1=3.2087029e-010             wkt1=3.857912e-008 pkt1=-3.319514e-015             kt2=-0.066969331               lkt2=3.0882088e-009 wkt2=2.0260742e-008             pkt2=-4.6329277e-015            ute=-2.0195803 lute=1.933839e-007              wute=1.0008578e-006             pute=-1.9916256e-013 ua1=2.5993531e-009             lua1=-1.9734905e-016            wua1=-1.0832502e-016 pua1=1.2514422e-022             ub1=-8.777109e-018             lub1=1.6721501e-024 wub1=5.0766552e-024             pub1=-1.2071184e-030            uc1=-1.9076744e-010 luc1=9.4252239e-017             wuc1=3.8850896e-016             puc1=-4.8067394e-023 at=309200.45                  lat=-0.059347591 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=-0.14900695                pat=2.597927e-008              vsat_ff=-13247.3 vsat_ss=364.054                    vsat_sf=-8487.14                   vsat_fs=14998.7 lvsat_ff=0.00229447                 lvsat_ss=0.00115062                 lvsat_sf=0.00152739 lvsat_fs=-0.00306155                wvsat_ff=0.0051026                  wvsat_ss=0.00629088 wvsat_sf=4e-09                      wvsat_fs=-0.0074791                 pvsat_ff=-1.04093e-09 pvsat_ss=-1.56139e-09               pvsat_sf=8e-16                      pvsat_fs=2.08186e-09 ags_ff=0.431863                   ags_ss=-0.305337                  ags_sf=-1.1264 ags_fs=0.374362                   lags_ff=-2.10862e-07               lags_ss=2.87232e-07 lags_sf=2.29785e-07                lags_fs=-7.63692e-08               wags_ff=-7.30438e-07 wags_ss=4.57832e-07                wags_sf=1.02052e-06                wags_fs=-4.2e-12 pags_ff=2.60231e-13                pags_ss=-2.60231e-13               pags_sf=-2.08185e-13 pags_fs=-2.3e-19                   at_ff=-28159.9                   at_sf=-16896 at_ss=28159.9                    at_fs=16896                      lat_ff=0.00574463 lat_sf=0.00344678                 lat_ss=-0.00574463                lat_fs=-0.00344678 wat_ff=0.0255129                  wat_sf=0.0153077                  wat_ss=-0.0255129 wat_fs=-0.0153077                 pat_ff=-5.20463e-09               pat_sf=-3.12278e-09 pat_ss=5.20463e-09                pat_fs=3.12278e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_12_mac.4 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=1.351e-06                  vth0=-0.51427127 lvth0=-4.4912792e-009            wvth0=-2.3959851e-008            pvth0=4.5480879e-015 k2=0.027258843                lk2=-6.8753191e-009            wk2=-2.1220692e-008 pk2=1.9826719e-015             cit=0.0012441903               lcit=3.4920343e-010 wcit=1.2596418e-010             pcit=-1.464941e-016             voff=-0.14346466 lvoff=-6.3359745e-009            wvoff=-1.9395282e-008            pvoff=3.3674775e-015 eta0=0.06679608                 weta0=3.0082752e-008             etab=-0.14741735 wetab=2.6505861e-008             u0=0.019946035                lu0=1.3665838e-009 wu0=4.6070809e-009             pu0=-1.1828646e-015            ua=1.258811e-009 lua=-1.2192925e-016            wua=-9.1599826e-016            pua=8.1488491e-023 ub=-2.055122e-019             lub=2.0218058e-025             wub=1.7708043e-024 pub=-2.3724708e-031            uc=-3.7714286e-011            luc=2.0771474e-017 wuc=3.9001143e-017             puc=-1.2411724e-023            vsat=72450.373 lvsat=-0.0011027087              wvsat=0.0018050833               pvsat=1.2648652e-009 a0=4.0046028                  la0=-9.5981131e-007            wa0=-1.6670576e-006 pa0=3.5822108e-013             ags=5.9116815                  lags=-4.6203218e-007 wags=-1.4266003e-006            pags=3.2405974e-013             keta=-0.10860686 lketa=2.2625349e-009             wketa=8.9156613e-008             pketa=-1.3342603e-014 pclm=0.63344537                 lpclm=-9.1772871e-009            wpclm=1.6039298e-007 ppclm=-1.8462599e-014            pdiblc2=0.0027536508               lpdiblc2=2.5425524e-010 wpdiblc2=1.6900495e-009             ppdiblc2=-3.447701e-016             agidl=1.2830406e-010 lagidl=-3.9994924e-018            wagidl=3.7660084e-017             pagidl=-1.1030982e-024 aigc=0.0068551817               laigc=-1.1961991e-011            waigc=-7.6369231e-011 paigc=-2.5946674e-018            aigsd=0.0059668795               laigsd=1.8027627e-011 waigsd=3.6488242e-011             paigsd=-3.1861963e-018            tvoff=0.000918222 ltvoff=-6.62503e-013              wtvoff=3.97058e-010               ptvoff=-5.09227e-018 kt1=-0.23183362                lkt1=-2.4010319e-009            wkt1=1.8156785e-008 pkt1=8.4664229e-016             kt2=-0.032414722               lkt2=-3.9609315e-009 wkt2=-1.006519e-008             pkt2=1.5535626e-015             ute=-1.0499167 lute=-4.4274761e-009            wute=-1.6672599e-007            pute=3.9024528e-014 ua1=6.9488612e-010             lua1=1.9116222e-016             wua1=1.5709784e-015 pua1=-2.1743367e-022            ub1=7.7992567e-019             lub1=-2.7748495e-025 wub1=-2.3413884e-024            pub1=3.0616253e-031             uc1=8.4238963e-011 luc1=3.8150931e-017             wuc1=3.2421197e-016             puc1=-3.4950807e-023 at=10812.968                  lat=0.0015234553 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=-0.033224207               pat=2.3595909e-009             letab=-4.3244943e-013 petab=6.5609751e-019             vsat_ff=-6963.39                   vsat_ss=15309.4 vsat_sf=-4413                      vsat_fs=1848.24                    lvsat_ff=0.00101253 lvsat_ss=-0.00189821                lvsat_sf=0.000696252                lvsat_fs=-0.000378856 wvsat_ff=0.00337514                 wvsat_ss=-0.00726938                wvsat_sf=0.00253132 wvsat_fs=0.00272604                 pvsat_ff=-6.88521e-10               pvsat_ss=1.20491e-09 pvsat_sf=-5.16389e-10               pvsat_fs=2e-15                      ags_ff=-0.974301 ags_ss=1.78526                    lags_ff=7.59954e-08                lags_ss=-1.39251e-07 wags_ff=8.82716e-07                wags_ss=-1.32407e-06               pags_ff=-6.88519e-14 pags_ss=1.03278e-13 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_12_mac.5 pmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=9e-007                     wmax=1.351e-06                  vth0=-0.59616193 lvth0=1.8961927e-009             wvth0=4.1813215e-008             pvth0=-5.822112e-016 k2=0.0039783965               lk2=-5.0594443e-009            wk2=1.1542835e-008 pk2=-5.7288321e-016            cit=0.0094033449               lcit=-2.8721063e-010 wcit=-5.2733318e-009            pcit=2.7465098e-016             voff=-0.20673273 lvoff=-1.4010648e-009            wvoff=2.3475884e-008             pvoff=2.3526537e-017 eta0=0.066797133                weta0=3.0081797e-008             etab=-0.32087101 wetab=6.5077776e-008             u0=0.035477085                lu0=1.5516191e-010 wu0=-8.3795638e-009            pu0=-1.6990633e-016            ua=2.5399611e-010 lua=-4.3553696e-017            wua=-8.8397341e-016            pua=7.8990552e-023 ub=3.0757673e-019             lub=1.6215964e-025             wub=9.5751219e-025 pub=-1.738103e-031             uc=1.2346667e-011             luc=1.686672e-017 wuc=6.552192e-017              puc=-1.4480344e-023            vsat=48802.426 lvsat=0.00074183115              wvsat=0.026342482                pvsat=-6.490519e-010 a0=-7.5648607                 la0=-5.7393159e-008            wa0=9.0205271e-006 pa0=-4.7541053e-013            ags=-2.7989296                 lags=2.1739548e-007 wags=6.5073486e-006             pags=-2.9478828e-013            keta=-0.11725185 lketa=2.9368444e-009             wketa=-1.0768649e-007            pketa=2.0111589e-015 pclm=0.2617378                  lpclm=1.9815903e-008             wpclm=1.8860407e-007 ppclm=-2.0663064e-014            pdiblc2=0.00032148148              lpdiblc2=4.4396444e-010 wpdiblc2=2.4267378e-009             ppdiblc2=-4.0223179e-016            agidl=-7.8456453e-011 lagidl=1.2127828e-017             wagidl=1.1657478e-016             pagidl=-7.2584442e-024 aigc=0.006857273                laigc=-1.2125114e-011            waigc=-2.8741157e-011 paigc=-6.3096572e-018            aigsd=0.0061646172               laigsd=2.6040867e-012 waigsd=5.8467506e-011             paigsd=-4.9005789e-018            tvoff=-0.000510203 ltvoff=1.10755e-010               wtvoff=1.87035e-009               ptvoff=-1.20009e-016 kt1=-0.32628496                lkt1=4.9661728e-009             wkt1=1.0982087e-007 pkt1=-6.3031563e-015            kt2=-0.14212147                lkt2=4.5961951e-009 wkt2=2.8462137e-008             pkt2=-1.451569e-015             ute=-1.118896 lute=9.5291271e-010             wute=2.3602148e-007             pute=7.6102254e-015 ua1=3.8440213e-009             lua1=-5.4470322e-017            wua1=-1.8692428e-015 pua1=5.0903579e-023             ub1=-2.9701376e-018            lub1=1.5019987e-026 wub1=1.6869879e-024             pub1=-8.050818e-033             uc1=5.7449965e-010 luc1=-8.9402338e-020            wuc1=-6.9080197e-017            puc1=-4.2740184e-024 at=53684.529                  lat=-0.0018205264 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=-0.036723864               pat=2.6325641e-009             letab=1.3528954e-008 petab=-3.0079533e-015            leta0=-8.2133422e-014            peta0=7.441288e-020 vsat_ff=17378.1                    vsat_ss=-26067.2                   vsat_sf=13033.6 vsat_fs=-8689.07                   lvsat_ff=-0.000886111               lvsat_ss=0.00132917 lvsat_sf=-0.000664584               lvsat_fs=0.000443056                wvsat_ff=-0.0157446 wvsat_ss=0.0236169                  wvsat_sf=-0.0118084                 wvsat_fs=0.0078723 pvsat_ff=8.02817e-10                pvsat_ss=-1.20423e-09               pvsat_sf=6.02113e-10 pvsat_fs=-4.01408e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_12_mac.6 pmos ( level=54                         lmin=9e-007                     lmax=9.023e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.52620375 lvth0=-1.0271625e-009            wvth0=5.8190815e-009             pvth0=1.5050565e-015 k2=0.019856783                lk2=-9.84774e-009              wk2=-1.9281855e-008 pk2=8.9179535e-015             cit=0.00087885845              lcit=1.1268006e-009 wcit=-4.8006604e-011            pcit=-2.3963797e-016            voff=-0.13309239 lvoff=-9.6398662e-009            wvoff=-1.5430919e-010            pvoff=2.4622233e-016 eta0=0.1                        etab=-0.15109442                wetab=2.9838581e-008 u0=0.012134061                lu0=2.6419234e-009             wu0=-8.2155302e-010 pu0=7.1489667e-016             ua=9.3046042e-010             lua=5.1073774e-017 wua=-2.9182404e-016            pua=2.9056765e-022             ub=8.7875458e-019 lub=1.7639822e-025             wub=-5.1925635e-026            pub=-1.0825168e-031 uc=-5.2922315e-011            luc=5.9970768e-017             wuc=-1.0294603e-016 puc=-1.0019385e-024            vsat=130796.57                  lvsat=-0.056142679 wvsat=-0.0030120476              pvsat=3.0653903e-008             a0=1.6667167 la0=-6.4646907e-007            wa0=-2.5694297e-008            pa0=3.908358e-013 ags=0.5899449                  lags=-1.2042422e-007            wags=-8.5039521e-008 pags=2.7384508e-013             keta=-0.011581329               lketa=1.1216984e-008 wketa=3.08628e-008               pketa=-3.0386629e-014            pclm=0.77591803 lpclm=1.4800767e-007             wpclm=1.6117154e-007             ppclm=-4.0619562e-013 pdiblc2=0.00055380988              lpdiblc2=-4.8364317e-010            wpdiblc2=-1.4310997e-010 ppdiblc2=1.2862724e-015             agidl=1.7205648e-010             lagidl=-6.9361575e-018 wagidl=-1.8000195e-017            pagidl=1.4607535e-023             aigc=0.0068018238 laigc=-3.3999986e-011            waigc=-2.5343698e-011            paigc=5.3538178e-018 aigsd=0.0060190044               laigsd=7.2898592e-011             waigsd=4.7133385e-011 paigsd=-6.4880623e-017            tvoff=0.00229365                 ltvoff=-1.48593e-009 wtvoff=-5.16288e-010              ptvoff=8.71036e-016               kt1=-0.19227935 lkt1=-3.898444e-008             wkt1=4.6721453e-009             pkt1=1.9362425e-014 kt2=-0.0474377                 lkt2=-1.7405205e-009            wkt2=-1.1273207e-008 pkt2=8.0550493e-015             ute=-0.97938499                lute=-7.0683177e-008 wute=2.3660964e-008             pute=5.7191733e-014             ua1=2.2538409e-009 lua1=2.6177702e-016             wua1=-1.1437311e-016            pua1=-9.7822737e-023 ub1=-2.6317584e-018            lub1=-3.4283107e-025            wub1=7.8063921e-026 pub1=2.1802493e-031             uc1=3.2287006e-010             luc1=-3.196532e-016 wuc1=1.1071235e-016             puc1=1.5849234e-022             at=128903.7 lat=0.0098535111               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              u0_ff=0.000199678 u0_ss=-0.000199678               u0_sf=0.000110932                u0_fs=-0.000110932 lu0_ff=-1.77313e-10               lu0_ss=1.77313e-10                lu0_sf=-9.85079e-11 lu0_fs=9.85079e-11                wu0_ff=-2e-16                     wu0_ss=2e-16 wu0_sf=-4.5e-16                   wu0_fs=4.5e-16                    pu0_ff=4e-22 pu0_ss=-4e-22                     pu0_sf=-2.2e-22                   pu0_fs=2.2e-22 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.7 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.52378198 lvth0=-3.177687e-009             wvth0=1.0126154e-008             pvth0=-2.3196241e-015 k2=0.009962078                lk2=-1.0612422e-009            wk2=-5.775859e-009 pk2=-3.0753707e-015            cit=0.002373555                lcit=-2.0048995e-010 wcit=-3.5533472e-010            pcit=3.3269397e-017             voff=-0.13020578 lvoff=-1.2203171e-008            wvoff=1.1129046e-009             pvoff=-8.7906355e-016 eta0=0.1                        etab=-0.15109442                wetab=2.9838581e-008 u0=0.010721391                lu0=3.8963745e-009             wu0=7.5092242e-010 pu0=-6.8146152e-016            ua=1.2213635e-009             lua=-2.0724815e-016 wua=-8.2527142e-017            pua=1.0471201e-022             ub=5.7586912e-019 lub=4.453605e-025              wub=1.5318172e-025             pub=-2.9038702e-031 uc=-2.5087662e-011            luc=3.5253596e-017             wuc=-9.3026936e-017 puc=-9.810089e-024             vsat=80512.667                  lvsat=-0.011490573 wvsat=0.032563367                pvsat=-9.3706541e-010            a0=1.0090829 la0=-6.2490285e-008            wa0=6.1746042e-007             pa0=-1.8028559e-013 ags=-0.041376927               lags=4.4018956e-007             wags=4.5690015e-007 pags=-2.0739735e-013            keta=0.032749059                lketa=-2.81484e-008 wketa=-2.8686882e-008            pketa=2.2493489e-014             pclm=1.1019734 lpclm=-1.4152952e-007            wpclm=-4.3642149e-007            ppclm=1.2446699e-013 pdiblc2=-0.00074111111             lpdiblc2=6.6624667e-010             wpdiblc2=9.7103067e-010 ppdiblc2=2.9691553e-016             agidl=1.9186716e-010             lagidl=-2.4528045e-017 wagidl=-3.7714648e-018            pagidl=1.9724229e-024             aigc=0.0067216027 laigc=3.7236362e-011             waigc=2.9343451e-011             paigc=-4.3208371e-017 aigsd=0.0062264338               laigsd=-1.1129871e-010            waigsd=-1.0704956e-010 paigsd=7.2033833e-017             tvoff=0.000119259                ltvoff=4.44922e-010 wtvoff=9.2651e-010                ptvoff=-4.10169e-016              kt1=-0.25083276 lkt1=1.301099e-008              wkt1=4.2634995e-008             pkt1=-1.4348585e-014 kt2=-0.060940876               lkt2=1.0250299e-008             wkt2=5.9650606e-009 pkt2=-7.2525327e-015            ute=-1.124714                  lute=5.8368994e-008 wute=1.5949782e-007             pute=-6.3431394e-014            ua1=2.3278537e-009 lua1=1.9605366e-016             wua1=-6.3110305e-017            pua1=-1.4334411e-022 ub1=-3.241586e-018             lub1=1.9869583e-025             wub1=2.9464452e-025 pub1=2.5701364e-032             uc1=-1.114144e-010             luc1=6.5991391e-017 wuc1=3.1242346e-016             puc1=-2.0627124e-023            at=213766.51 lat=-0.065504662               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=-0.0092519848 pat=8.2157625e-009             vsat_ff=3390.47                    vsat_ss=-4363.74 vsat_sf=7819.13                    vsat_fs=-12247.8                   lvsat_ff=-0.00301069 lvsat_ss=0.003875                   lvsat_sf=-0.00694334                lvsat_fs=0.010876 wvsat_ff=0.00133745                 wvsat_ss=-0.00133746                wvsat_sf=-0.00267492 wvsat_fs=0.00668729                 pvsat_ff=-1.18766e-09               pvsat_ss=1.18766e-09 pvsat_sf=2.37532e-09                pvsat_fs=-5.93831e-09               ags_ff=0.194667 ags_ss=-0.194667                  ags_fs=-0.489911                  ags_sf=-0.295244 lags_ff=-1.72864e-07               lags_ss=1.72864e-07                lags_fs=4.35041e-07 lags_sf=2.62177e-07                wags_ff=4.7e-13                    wags_ss=-4.7e-13 wags_fs=2.67491e-07                wags_sf=2.67491e-07                pags_ff=-4.2e-19 pags_ss=4.2e-19                    pags_fs=-2.37532e-13               pags_sf=-2.37532e-13 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.8 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.51961828 lvth0=-5.0013903e-009            wvth0=4.2946009e-009             pvth0=2.3459629e-016 k2=0.02410858                 lk2=-7.2574099e-009            wk2=-1.78943e-008 pk2=2.2325064e-015             cit=0.0012225611               lcit=3.0364534e-010 wcit=-2.0018382e-010            pcit=-3.4686697e-017            voff=-0.13608182 lvoff=-9.6294673e-009            wvoff=-6.0761984e-009            pvoff=2.2697636e-015 eta0=0.1                        etab=-0.15109442                wetab=2.9838581e-008 u0=0.016239163                lu0=1.4795903e-009             wu0=-2.958429e-009 pu0=9.432344e-016              ua=1.3777043e-009             lua=-2.7572544e-016 wua=2.4177469e-016             pua=-3.7332195e-023            ub=1.7770942e-018 lub=-8.0776061e-026            wub=-1.0137432e-024            pub=2.2072609e-031 uc=3.514203e-011              luc=8.8729909e-018             wuc=-1.8553345e-016 puc=3.0707763e-023             vsat=35991.529                  lvsat=0.0080096858 wvsat=0.056452766                pvsat=-1.1400622e-008            a0=2.6730206 la0=-7.9129498e-007            wa0=-9.1503469e-008            pa0=1.3024059e-013 ags=-2.2540966                 lags=1.4093608e-006             wags=6.236833e-007 pags=-2.8044836e-013            keta=0.018107297                lketa=-2.1735309e-008 wketa=2.8893416e-008             pketa=-2.7266815e-015            pclm=0.87017009 lpclm=-3.9999657e-008            wpclm=-2.7827287e-007            ppclm=5.5197893e-014 pdiblc2=-0.0013660684              lpdiblc2=9.3997795e-010             wpdiblc2=2.4874733e-009 ppdiblc2=-3.6728636e-016            agidl=1.3106828e-010             lagidl=2.1018642e-018 wagidl=-9.4151222e-019            pagidl=7.3290367e-025             aigc=0.006807923 laigc=-5.7193738e-013            waigc=-4.5286743e-011            paigc=-1.0520346e-017 aigsd=0.0058851095               laigsd=3.8201328e-011             waigsd=1.0279076e-010 paigsd=-1.9876226e-017            tvoff=0.00133927                 ltvoff=-8.94426e-011 wtvoff=-3.54187e-010              ptvoff=1.50777e-016               kt1=-0.1953596 lkt1=-1.1286255e-008            wkt1=-6.554793e-009             pkt1=7.1965418e-015 kt2=-0.037172139               lkt2=-1.604078e-010             wkt2=-6.735514e-009 pkt2=-1.689681e-015             ute=-0.88702626                lute=-4.5738243e-008 wute=-2.5236201e-008            pute=1.7482107e-014             ua1=3.0364834e-009 lua1=-1.1432614e-016            wua1=-5.0436505e-016            pua1=4.9925471e-023 ub1=-3.4489545e-018            lub1=2.8952323e-025             wub1=2.4934713e-025 pub1=4.554162e-032              uc1=9.7124287e-011             luc1=-2.5348555e-017 wuc1=1.2767905e-016             puc1=6.0290924e-023             at=119744.2 lat=-0.024322888               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=0.022640421 pat=-5.7531114e-009            vsat_ff=-4776.47                   vsat_ss=3807.68 vsat_sf=-16809.4                   vsat_fs=16971.4                    lvsat_ff=0.00056641 lvsat_ss=0.000295933                lvsat_sf=0.00384392                 lvsat_fs=-0.00192196 wvsat_ff=-0.002572                  wvsat_ss=0.00317103                 wvsat_sf=0.0075399 wvsat_fs=-0.00926637                pvsat_ff=5.24699e-10                pvsat_ss=-7.87044e-10 pvsat_sf=-2.09878e-09               pvsat_fs=1.04939e-09                ags_ff=-0.374359 ags_ss=-0.0644438                 ags_fs=0.942137                   ags_sf=0.567778 lags_ff=7.63693e-08                lags_ss=1.15827e-07                lags_fs=-1.92196e-07 lags_sf=-1.15827e-07               wags_ff=3.3e-13                    wags_ss=2.39587e-07 wags_fs=-5.14407e-07               wags_sf=-5.14407e-07               pags_ff=-4e-20 pags_ss=-1.04939e-13               pags_fs=1.04939e-13                pags_sf=1.04939e-13 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.9 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.54932553 lvth0=1.0588895e-009             wvth0=7.7993127e-009             pvth0=-4.8036492e-016 k2=0.01414577                 lk2=-5.2249968e-009            wk2=-9.3402485e-009 pk2=4.8747995e-016             cit=0.0018553249               lcit=1.7456154e-010 wcit=-4.2772375e-010            pcit=1.1731449e-017             voff=-0.17301288 lvoff=-2.0955305e-009            wvoff=7.3754113e-009             pvoff=-4.743648e-016 eta0=0.1                        etab=-0.15109801                wetab=2.9840546e-008 u0=0.023283481                lu0=4.254945e-011              wu0=1.5833548e-009 pu0=1.6710515e-017             ua=-1.6982755e-010            lua=3.9971061e-017 wua=3.7834822e-016             pua=-6.5193194e-023            ub=2.1313316e-018 lub=-1.5304051e-025            wub=-3.4637622e-025            pub=8.4583229e-032 uc=1.0168861e-010             luc=-4.7025117e-018            wuc=-8.7297882e-017 puc=1.0667708e-023             vsat=83832.676                  lvsat=-0.0017499081 wvsat=-0.0085072833              pvsat=1.8512279e-009             a0=2.0320144 la0=-6.6052972e-007            wa0=1.2010748e-007             pa0=8.7071959e-014 ags=6.8301143                  lags=-4.4381825e-007            wags=-2.2587004e-006 pags=3.0755791e-013             keta=-0.037947778               lketa=-1.0300073e-008 wketa=2.5139487e-008             pketa=-1.96088e-015              pclm=0.81337358 lpclm=-2.841317e-008             wpclm=-2.6219733e-009            ppclm=-1.0348893e-015 pdiblc2=0.0033912698               lpdiblc2=-3.0519048e-011            wpdiblc2=1.1123667e-009 ppdiblc2=-8.67646e-017              agidl=1.7309033e-010             lagidl=-6.4706337e-018 wagidl=-2.9162772e-018            pagidl=1.1357557e-024             aigc=0.0068432804 laigc=-7.7848401e-012            waigc=-6.5586645e-011            paigc=-6.3791659e-018 aigsd=0.0059942673               laigsd=1.5933138e-011             waigsd=1.1674891e-011 paigsd=-1.2885897e-018            tvoff=0.000668911                ltvoff=4.73106e-011 wtvoff=6.22934e-010               ptvoff=-4.85559e-017              kt1=-0.25588901 lkt1=1.0617445e-009             wkt1=3.9950966e-008             pkt1=-2.2906332e-015 kt2=-0.0074151625              lkt2=-6.2308309e-009            wkt2=-3.2714791e-008 pkt2=3.6100915e-015             ute=-1.3589699                 lute=5.0538259e-008 wute=1.1327622e-007             pute=-1.0774428e-014            ua1=2.6187934e-009 lua1=-2.9117379e-017            wua1=-1.7208159e-016            pua1=-1.7860354e-023 ub1=-2.2387569e-018            lub1=4.2642939e-026             wub1=3.9353809e-025 pub1=1.6126664e-032             uc1=-3.4003932e-010            luc1=6.3832822e-017 wuc1=7.0860809e-016             puc1=-5.82186e-023              at=-17045.157 lat=0.0035821398               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=-0.0079847459 pat=4.9442272e-010             letab=7.34162e-013               petab=-4.0085245e-019 vsat_ff=-4176.99                   vsat_ss=10391.3                    vsat_sf=2353.18 vsat_fs=12223.8                    lvsat_ff=0.000444104                lvsat_ss=-0.00104713 lvsat_sf=-6.5248e-05                lvsat_fs=-0.000953457               wvsat_ff=0.000850633 wvsat_ss=-0.00281367                wvsat_sf=-0.00359884                wvsat_fs=-0.0066742 pvsat_ff=-1.73529e-10               pvsat_ss=4.33823e-10                pvsat_sf=1.7353e-10 pvsat_fs=5.20588e-10                ags_ss=0.814921                   lags_ss=-6.35638e-08 wags_ss=-4.44947e-07               pags_ss=3.47058e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.10 pmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.5474461 lvth0=9.1229362e-010             wvth0=-2.3233323e-009            pvth0=3.0920138e-016 k2=0.030217995                lk2=-6.4786304e-009            wk2=-1.2230242e-008 pk2=7.128994e-016              cit=0.0034878125               lcit=4.7227502e-011 wcit=8.6140566e-011             pcit=-2.8349968e-017            voff=-0.18055851 lvoff=-1.5069717e-009            wvoff=-2.3795946e-010            pvoff=1.1947812e-016 eta0=0.1                        etab=-0.33438299                wetab=7.7319626e-008 u0=0.024049126                lu0=-1.7170831e-011            wu0=1.9741673e-009 pu0=-1.3772865e-017            ua=1.6713812e-010             lua=1.3687739e-017 wua=-8.0528006e-016            pua=2.7129812e-023             ub=1.1110998e-019 lub=4.5367784e-027             wub=1.1355111e-024             pub=-3.100398e-032 uc=-9.5985185e-011            luc=1.0716044e-017             wuc=1.6367058e-016 puc=-8.9078323e-024            vsat=44595.734                  lvsat=0.0013105734 wvsat=0.030153746                pvsat=-1.1643324e-009            a0=0.54030873 la0=-5.4417668e-007            wa0=1.6772436e-006             pa0=-3.438466e-014 ags=-0.5696224                 lags=1.3336122e-007             wags=4.4875962e-006 pags=-2.1865323e-013            keta=-0.26475926                lketa=7.3912222e-009 wketa=2.5955222e-008             pketa=-2.0245073e-015            pclm=0.4883107 lpclm=-3.0582652e-009            wpclm=-1.6670974e-008            ppclm=6.0932812e-017 pdiblc2=0.0058648148               lpdiblc2=-2.2345556e-010            wpdiblc2=-2.5955222e-009 ppdiblc2=2.0245073e-016             agidl=8.6263082e-011             lagidl=3.0189173e-019 wagidl=-3.2661122e-017            pagidl=3.4558537e-024             aigc=0.0071779899 laigc=-3.389218e-011             waigc=-3.1931062e-010            paigc=1.3411304e-017 aigsd=0.0061306372               laigsd=5.2962861e-012             waigsd=8.9253378e-011 paigsd=-7.3397116e-018            tvoff=0.0020942                  ltvoff=-6.38622e-011 wtvoff=-4.89239e-010              ptvoff=3.81936e-017               kt1=-0.18306268 lkt1=-4.6187089e-009            wkt1=-1.9938517e-008            pkt1=2.3807465e-015 kt2=-0.15397088                lkt2=5.2005146e-009             wkt2=3.9197696e-008 pkt2=-1.9990825e-015            ute=-0.77912567                lute=5.310409e-009 wute=-7.1810466e-008            pute=3.6623338e-015             ua1=3.1970113e-009 lua1=-7.4218379e-017            wua1=-1.2830518e-015            pua1=6.8795318e-023 ub1=-3.1896204e-018            lub1=1.1681029e-025             wub1=1.8858393e-024 pub1=-1.0027283e-031            uc1=8.1926869e-010             luc1=-2.6593204e-017 wuc1=-2.9084095e-016            puc1=1.9738425e-023             at=7295.1289 lat=0.0016835976               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=0.0053049323 pat=-5.4217217e-010            letab=1.4296962e-008             petab=-3.7037691e-015 u0_ff=0.00128844                 u0_ss=-0.00229055                u0_fs=-0.00114528 lu0_ff=-1.00498e-10               lu0_ss=1.78663e-10                lu0_fs=8.93316e-11 wu0_ff=-1.16732e-09               wu0_ss=2.07524e-09                wu0_fs=1.03762e-09 pu0_ff=9.10512e-17                pu0_ss=-1.61869e-16               pu0_fs=-8.09344e-17 vsat_ff=5238.82                    vsat_ss=-13054.5                   vsat_sf=4379.86 lvsat_ff=-0.000290328               lvsat_ss=0.000781652                lvsat_sf=-0.000223329 wvsat_ff=-0.00474637                wvsat_ss=0.0118274                  wvsat_sf=-0.00396815 pvsat_ff=2.63037e-10                pvsat_ss=-7.08176e-10               pvsat_sf=2.02336e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.11 pmos ( level=54                         lmin=9e-007                     lmax=9.023e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.51143929 lvth0=-3.0173825e-009            wvth0=-2.2423108e-009            pvth0=2.5917167e-015 k2=-0.017915255               lk2=1.2221094e-008             wk2=1.3416776e-009 pk2=-3.13163e-015              cit=0.00058409469              lcit=1.0665578e-009 wcit=1.1293441e-010             pcit=-2.0674545e-016            voff=-0.13040638 lvoff=-8.5834378e-009            wvoff=-1.62087e-009              pvoff=-3.3058758e-016 eta0=0.1                        etab=-0.1379094                 wetab=2.2639562e-008 u0=0.0097552428               lu0=4.0076638e-009             wu0=4.7728172e-010 pu0=-3.0797609e-017            ua=4.7432303e-010             lua=4.9544608e-016 wua=-4.2773024e-017            pua=4.7940372e-023             ub=7.1872339e-019 lub=-9.7477098e-027            wub=3.5451395e-026             pub=-6.6160083e-033 uc=-2.9024254e-010            luc=1.0144737e-016             wuc=2.6630815e-017 puc=-2.3648164e-023            vsat=122299.52                  lvsat=0.025594167 wvsat=0.0016273432               pvsat=-1.3974415e-008            a0=1.5759176 la0=-3.7845296e-008            wa0=2.3881997e-008             pa0=5.8527215e-014 ags=0.30027603                 lags=2.7918763e-007             wags=7.3119682e-008 pags=5.5657012e-014             keta=0.078740387                lketa=-7.2566599e-008 wketa=-1.8452857e-008            pketa=1.5359207e-014             pclm=1.2191145 lpclm=-9.6338435e-007            wpclm=-8.0813738e-008            ppclm=2.0062442e-013 pdiblc2=0.00017963786              lpdiblc2=2.8794149e-009             wpdiblc2=6.1187951e-011 ppdiblc2=-5.499573e-016             agidl=1.2025889e-010             lagidl=5.6856076e-017 wagidl=1.0281285e-017             pagidl=-2.0223024e-023            aigc=0.0067953326 laigc=5.2928514e-012             waigc=-2.1799482e-011            paigc=-1.6100072e-017 aigsd=0.0061041973               laigsd=-1.0266085e-010            waigsd=6.1805597e-013 paigsd=3.0974833e-017             tvoff=0.00126248                 ltvoff=-1.8309e-010 wtvoff=4.6731e-011                ptvoff=1.59683e-016               kt1=-0.19693793 lkt1=-1.1758836e-008            wkt1=7.215729e-009              pkt1=4.4972456e-015 kt2=-0.084526637               lkt2=2.6313797e-008             wkt2=8.9773517e-009 pkt2=-7.2626079e-015            ute=-0.93671255                lute=2.4676038e-008 wute=3.6181097e-010             pute=5.125602e-015              ua1=2.2236367e-009 lua1=3.102397e-017              wua1=-9.7881602e-017            pua1=2.8168428e-023 ub1=-2.7976507e-018            lub1=2.5111763e-025             wub1=1.6864116e-025 pub1=-1.0627105e-031            uc1=6.6525557e-010             luc1=-2.4390398e-016 wuc1=-7.6230139e-017            puc1=1.1713326e-022             at=125582.07 lat=0.039708336                jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=0.0018136109 pat=-1.6300734e-008            u0_ff=0.000199677                u0_ss=-0.000199677 u0_sf=0.000110932                u0_fs=-0.000110932               lu0_ff=-1.77313e-10 lu0_ss=1.77313e-10                lu0_sf=-9.85074e-11               lu0_fs=9.85074e-11 wu0_ff=-3.5e-16                   wu0_ss=3.5e-16                    wu0_sf=3e-18 wu0_fs=-3e-18                     pu0_ff=-2.1e-23                   pu0_ss=2.1e-23 pu0_sf=-4.5e-23                   pu0_fs=4.5e-23                    ags_ff=0.0340191 ags_ss=-0.0340191                 lags_ff=-3.0209e-08                lags_ss=3.0209e-08 wags_ff=-1.85744e-08               wags_ss=1.85744e-08                pags_ff=1.64941e-14 pags_ss=-1.64941e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.12 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.49897398 lvth0=-1.4086581e-008            wvth0=-3.4190173e-009            pvth0=3.6366321e-015 k2=0.0035517881               lk2=-6.8416396e-009            wk2=-2.2758407e-009 pk2=8.0726255e-017             cit=0.0018892653               lcit=-9.2433619e-011 wcit=-9.0912536e-011            pcit=-2.5729359e-017            voff=-0.1171015 lvoff=-2.0398172e-008            wvoff=-6.0420352e-009            pvoff=3.5954071e-015 eta0=0.1                        etab=-0.1379094                 wetab=2.2639562e-008 u0=0.0099488542               lu0=3.8357369e-009             wu0=1.1727274e-009 pu0=-6.483534e-016             ua=9.0063152e-010             lua=1.1688414e-016 wua=9.2592509e-017             pua=-7.2264221e-023            ub=8.75709e-019 lub=-1.4915093e-025            wub=-1.0530848e-026            pub=3.4216223e-032 uc=-1.9148681e-010            luc=1.3752292e-017             wuc=-2.1729991e-018 puc=1.9296232e-024             vsat=161298.09                  lvsat=-0.0090365616 wvsat=-0.011545472               pvsat=-2.2769554e-009            a0=1.9385962 la0=-3.599039e-007             wa0=1.0994616e-007             pa0=-1.7897757e-014 ags=0.88358841                 lags=-2.3879376e-007            wags=-4.8130917e-008 pags=1.6332754e-013             keta=-0.03551067                lketa=2.888834e-008 wketa=8.5829297e-009             pketa=-8.6485712e-015            pclm=-0.20861623 lpclm=3.0444055e-007             wpclm=2.7916046e-007             ppclm=-1.1903267e-013 pdiblc2=0.0024575407               lpdiblc2=8.5663716e-010             wpdiblc2=-7.7543324e-010 ppdiblc2=1.9296232e-016             agidl=2.146799e-010              lagidl=-2.698978e-017 wagidl=-1.6227222e-017            pagidl=3.3165303e-024             aigc=0.0068606019 laigc=-5.2666306e-011            waigc=-4.6550109e-011            paigc=5.8784862e-018 aigsd=0.0059345251               laigsd=4.8007987e-011             waigsd=5.2332534e-011 paigsd=-1.4947624e-017            tvoff=0.00155908                 ltvoff=-4.46475e-010 wtvoff=1.40368e-010               ptvoff=7.65338e-017               kt1=-0.19331564 lkt1=-1.4975427e-008            wkt1=1.1230647e-008             pkt1=9.3199836e-016 kt2=-0.059864437               lkt2=4.4137636e-009             wkt2=5.3773252e-009 pkt2=-4.0657844e-015            ute=-0.83230602                lute=-6.8036965e-008 wute=-1.5694709e-010            pute=5.5862592e-015             ua1=2.1422506e-009 lua1=1.0329485e-016             wua1=3.8229011e-017             pua1=-9.2697797e-023 ub1=-2.7450647e-018            lub1=2.0442124e-025             wub1=2.3543922e-026 pub1=2.2575289e-032             uc1=2.9862501e-010             luc1=8.1663953e-017 wuc1=8.8541938e-017             puc1=-2.9184344e-023            at=231255.6 lat=-0.054129757               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=-0.018801027 pat=2.0050644e-009             vsat_ff=9819.87                    vsat_ss=-11788.2 vsat_sf=5904.89                    lvsat_ff=-0.00872005                lvsat_ss=0.0104678 lvsat_sf=-0.00524354                wvsat_ff=-0.002173                  wvsat_ss=0.00271625 wvsat_sf=-0.00162975                pvsat_ff=1.92962e-09                pvsat_ss=-2.41203e-09 pvsat_sf=1.44722e-09                ags_ff=0.194666                   ags_ss=-0.194666 ags_sf=0.393659                   lags_ff=-1.72864e-07               lags_ss=1.72864e-07 lags_sf=-3.49569e-07               wags_ff=-4e-14                     wags_ss=4e-14 wags_sf=-1.0865e-07                pags_ff=3.9e-20                    pags_ss=-3.9e-20 pags_sf=9.64812e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.13 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.51948706 lvth0=-5.1018518e-009            wvth0=4.2229548e-009             pvth0=2.8944825e-016 k2=-0.007218623               lk2=-2.1241995e-009            wk2=-7.8964726e-010 pk2=-5.7022647e-016            cit=0.00084727984              lcit=3.6395599e-010 wcit=4.7197691e-012             pcit=-6.7616309e-017            voff=-0.14945733 lvoff=-6.226319e-009             wvoff=1.226829e-009              pvoff=4.1164462e-016 eta0=0.1                        etab=-0.1379094                 wetab=2.2639562e-008 u0=0.0095143687               lu0=4.0260416e-009             wu0=7.1330871e-010 pu0=-4.47128e-016              ua=2.0937856e-009             lua=-4.0571737e-016 wua=-1.492057e-016             pua=3.3643394e-023             ub=-5.8431271e-019 lub=4.9033857e-025             wub=2.7558496e-025             pub=-9.11025e-032 uc=-3.7393085e-010            luc=9.366278e-017              wuc=3.7820345e-017 puc=-1.5587462e-023            vsat=202797.67                  lvsat=-0.027213379 wvsat=-0.034623387               pvsat=7.8311715e-009             a0=2.6440423 la0=-6.688893e-007             wa0=-7.5681357e-008            pa0=6.3407093e-014 ags=-1.4933081                 lags=8.0228689e-007             wags=2.0829276e-007 pags=5.1013973e-014             keta=0.14898875                 lketa=-5.1922405e-008 wketa=-4.2567856e-008            pketa=1.3755473e-014             pclm=0.32624489 lpclm=7.0171375e-008             wpclm=1.8710289e-008             ppclm=-4.955491e-015 pdiblc2=0.0047833618               lpdiblc2=-1.6207248e-010            wpdiblc2=-8.7011556e-010 ppdiblc2=2.3443317e-016             agidl=1.5223605e-010             lagidl=3.6062904e-019 wagidl=-1.2499112e-017            pagidl=1.6836181e-024             aigc=0.0067558394 laigc=-6.7803327e-012            waigc=-1.6849086e-011            paigc=-7.130562e-018 aigsd=0.0060627953               laigsd=-8.174353e-012             waigsd=5.77427e-012 paigsd=5.4448959e-018             tvoff=-0.000322309               ltvoff=3.77574e-010 wtvoff=5.53035e-010               ptvoff=-1.04214e-016              kt1=-0.2408573 lkt1=5.847821e-009              wkt1=1.8286953e-008             pkt1=-2.1586639e-015 kt2=-0.038179844               lkt2=-5.0840881e-009            wkt2=-6.1853068e-009 pkt2=9.9864845e-016             ute=-0.85341479                lute=-5.8791325e-008 wute=-4.3588067e-008            pute=2.460909e-014              ua1=2.6528625e-009 lua1=-1.2035318e-016            wua1=-2.9490804e-016            pua1=5.321623e-023 ub1=-3.0674015e-018            lub1=3.4560475e-025             wub1=4.1019206e-026 pub1=1.4921115e-032             uc1=3.1823522e-010             luc1=7.3074682e-017 wuc1=6.9524838e-018             puc1=6.5518373e-024             at=196309.22 lat=-0.038823242               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=-0.019164081 pat=2.1640817e-009             vsat_ff=-18031.9                   vsat_ss=20964.6 vsat_sf=-6066.67                   lvsat_ff=0.00347904                 lvsat_ss=-0.00387786 lvsat_sf=3.3e-09                    wvsat_ff=0.00466542                 wvsat_ss=-0.00619672 wvsat_sf=0.0016744                  pvsat_ff=-1.06561e-09               pvsat_ss=1.49185e-09 pvsat_sf=-2e-16                     ags_ff=-0.374359                  ags_ss=0.374359 ags_sf=-0.757037                  lags_ff=7.63697e-08                lags_ss=-7.63697e-08 lags_sf=1.54436e-07                wags_ff=-2.2e-13                   wags_ss=2.2e-13 wags_sf=2.08942e-07                pags_ff=1.3e-20                    pags_ss=-1.3e-20 pags_sf=-4.26242e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.14 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.55059797 lvth0=1.2447737e-009             wvth0=8.4940624e-009             pvth0=-5.818577e-016 k2=0.0069324468               lk2=-5.0110178e-009            wk2=-5.401774e-009 pk2=3.7064738e-016             cit=0.0016846486               lcit=1.9313277e-010 wcit=-3.3453447e-010            pcit=1.5915559e-018             voff=-0.16708502 lvoff=-2.6302698e-009            wvoff=4.1387984e-009             pvoff=-1.8239714e-016 eta0=0.1                        etab=-0.13790941                wetab=2.2639569e-008 u0=0.031002122                lu0=-3.5746019e-010            wu0=-2.6310235e-009 pu0=2.3511578e-016             ua=5.3464614e-10              lua=-8.7652908e-17 wua=-6.2944194e-18             pua=4.4894929e-24              ub=1.9719038e-018 lub=-3.1129591e-026            wub=-2.593286e-025             pub=1.8019866e-032 uc=4.1041953e-011             luc=9.0083276e-018             wuc=-5.4184807e-017 puc=3.1815893e-024             vsat=59299.353                  lvsat=0.0020602772 wvsat=0.0048879112               pvsat=-2.2913332e-010            a0=1.7770987 la0=-4.920328e-007             wa0=2.5929144e-007             pa0=-4.9273582e-015 ags=0.55892505                 lags=3.8363133e-007             wags=1.1653689e-006 pags=-1.4422956e-013            keta=-0.10359286                lketa=-3.9575698e-010 wketa=6.0981701e-008             pketa=-7.3686367e-015            pclm=0.83144973 lpclm=-3.2890413e-008            wpclm=-1.2491556e-008            ppclm=1.4096853e-015 pdiblc2=0.0046010582               lpdiblc2=-1.2488254e-010            wpdiblc2=4.5182222e-010 ppdiblc2=-3.5242133e-017            agidl=1.9825666e-010             lagidl=-9.027576e-018 wagidl=-1.6657094e-017            pagidl=2.5318462e-024             aigc=0.0068042148 laigc=-1.6648911e-011            waigc=-4.4256824e-011            paigc=-1.5393834e-018 aigsd=0.0059046186               laigsd=2.4093698e-011             waigsd=6.0623052e-011 paigsd=-5.7442556e-018            tvoff=0.00153426                 ltvoff=-1.16588e-012 wtvoff=1.50453e-010               ptvoff=-2.20878e-017              kt1=-0.21029887 lkt1=-3.860993e-010             wkt1=1.505875e-008              pkt1=-1.5001104e-015 kt2=-0.065096413               lkt2=4.0689185e-010             wkt2=-1.2208284e-009 pkt2=-1.4105149e-017            ute=-1.4111464                 lute=5.4985935e-008 wute=1.4176462e-007             pute=-1.3202859e-014            ua1=2.7384776e-009 lua1=-1.3781865e-016            wua1=-2.3742916e-016            pua1=4.149054e-023 ub1=-2.3231324e-018            lub1=1.9377384e-025             wub1=4.3960707e-025 pub1=-6.6390809e-032            uc1=8.4475831e-010             luc1=-3.4336029e-017 wuc1=6.1708584e-017             puc1=-4.6184072e-024            at=-4076.1793 lat=0.0020553792               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=-0.015065808 pat=1.328034e-009              letab=2.2978387e-015             petab=-1.2546199e-021 vsat_ff=301.579                    vsat_ss=1928.04                    vsat_sf=-8570.37 lvsat_ff=-0.00026099                lvsat_ss=5.61338e-06                lvsat_sf=0.000510755 wvsat_ff=-0.00159466                wvsat_ss=0.00180729                 wvsat_sf=0.00236542 pvsat_ff=2.11453e-10                pvsat_ss=-1.40969e-10               pvsat_sf=-1.40969e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.15 pmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.54918675 lvth0=1.1346988e-009             wvth0=-1.3729356e-009            pvth0=1.8776815e-016 k2=0.011413998                lk2=-5.3605787e-009            wk2=-1.9632588e-009 pk2=1.024432e-016              cit=0.0046431006               lcit=-3.7626487e-011 wcit=-5.446467e-010             pcit=1.798031e-017              voff=-0.17847547 lvoff=-1.7418149e-009            wvoff=-1.3752998e-009            pvoff=2.4770252e-016 eta0=0.1                        etab=-0.29022609                wetab=5.3209961e-008 u0=0.02241804                 lu0=3.1209828e-010             wu0=2.8647403e-009 pu0=-1.935538e-016             ua=-2.1529382e-09             lua=1.2197867e-16 wua=4.6148162e-16              pua=-3.1997039e-23             ub=2.7703957e-018 lub=-9.3411964e-026            wub=-3.1645896e-025            pub=2.2476034e-032 uc=1.858321e-010              luc=-2.2853037e-018            wuc=9.7983407e-018 puc=-1.8090962e-024            vsat=98352.665                  lvsat=-0.00098588106 wvsat=0.00080246137              pvsat=8.9531765e-011             a0=3.0209312 la0=-5.8905174e-007            wa0=3.2282376e-007             pa0=-9.8828786e-015 ags=12.402157                  lags=-5.4014076e-007            wags=-2.5949953e-006 pags=1.4907885e-013             keta=-0.049691358               lketa=-4.6000741e-009 wketa=-9.1471852e-008            pketa=4.5227404e-015             pclm=0.38962963 lpclm=1.5715556e-009             wpclm=3.7208889e-008             ppclm=-2.4669493e-015 pdiblc2=-0.00081975309             lpdiblc2=2.9794074e-010             wpdiblc2=1.0542519e-009 ppdiblc2=-8.2231644e-017            agidl=1.4898806e-011             lagidl=5.2743366e-018 wagidl=6.3037721e-018             pagidl=7.4089873e-025             aigc=0.0066955956 laigc=-8.1766174e-012            waigc=-5.5923371e-011            paigc=-6.2939278e-019 aigsd=0.0062377865               laigsd=-1.8933975e-012            waigsd=3.0749831e-011 paigsd=-3.4141444e-018            tvoff=0.0024066                  ltvoff=-6.9208e-011 wtvoff=-6.59805e-010              ptvoff=4.11124e-017               kt1=-0.19535009 lkt1=-1.5521039e-009            wkt1=-1.3229591e-008            pkt1=7.0638019e-016 kt2=-0.074764013               lkt2=1.1609646e-009             wkt2=-4.0492505e-009 pkt2=2.0651177e-016             ute=-0.8134008                 lute=8.3617743e-009 wute=-5.3096241e-008            pute=1.9962883e-015             ua1=-2.7202452e-010 lua1=9.7000513e-017             wua1=6.1104182e-016             pua1=-2.4690197e-023 ub1=1.497659e-018              lub1=-1.0424788e-025            wub1=-6.7341521e-025 pub1=2.0424929e-032             uc1=2.347575e-010              luc1=1.3244034e-017 wuc1=2.8302162e-017             puc1=-2.0127063e-024            at=-3631.6815 lat=0.0020207084               jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)' jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)'                              wat=0.011270971 pat=-7.262347e-010             letab=1.1880703e-008             petab=-2.3844919e-015 u0_ff=-0.00171792                u0_ss=0.00305407                 u0_fs=0.00152704 lu0_ff=1.33997e-10                lu0_ss=-2.38218e-10               lu0_fs=-1.19109e-10 wu0_ff=4.74145e-10                wu0_ss=-8.42924e-10               wu0_fs=-4.21462e-10 pu0_ff=-3.69833e-17               pu0_ss=6.57481e-17                pu0_fs=3.2874e-17 vsat_ff=-6077.54                   vsat_ss=7642.51                    vsat_sf=-5839.81 vsat_mc=-1543.82                   lvsat_ff=0.000236581                lvsat_ss=-0.000440114 lvsat_sf=0.000297772                lvsat_mc=0.000120418                wvsat_ff=0.00143237 wvsat_ss=0.000526826                wvsat_sf=0.00161179                 wvsat_mc=0.000842924 pvsat_ff=-2.46552e-11               pvsat_ss=-4.10922e-11               pvsat_sf=-8.21851e-11 pvsat_mc=-6.57481e-11 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.16 pmos ( level=54                         lmin=9e-007                     lmax=9.023e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.52322044 lvth0=9.9906703e-009             wvth0=1.0092856e-009             pvth0=-9.9850591e-016 k2=-0.028122554               lk2=3.2161764e-009             wk2=4.1588921e-009 pk2=-6.4627263e-016            cit=0.0013601566               lcit=3.0669783e-010 wcit=-1.0125868e-010            pcit=2.9759136e-018             voff=-0.1452081 lvoff=-6.1509176e-009            wvoff=2.4644034e-009             pvoff=-1.0019631e-015 eta0=0.11407407                 weta0=-3.8844444e-009            etab=-0.063634 wetab=2.139552e-009              u0=0.010908525                lu0=4.2219741e-009 wu0=1.5897592e-010             pu0=-8.9947229e-017            ua=3.526916e-010 lua=5.5535708e-016             wua=-9.2027494e-018            pua=3.1404935e-023 ub=9.5465249e-019             lub=1.6627774e-025             wub=-2.9665037e-026 pub=-5.5199033e-032            uc=-2.7000786e-010            luc=5.0828534e-017 wuc=2.1046045e-017             puc=-9.6773649e-024            vsat=121793.49 lvsat=-0.024039283               wvsat=0.0017670079               pvsat=-2.75583e-010 a0=1.4144165                  la0=3.8072501e-007             wa0=6.8456294e-008 pa0=-5.6998189e-014            ags=0.43002277                 lags=6.1506205e-007 wags=3.7309581e-008             pags=-3.7044327e-014            keta=0.03048152 lketa=-2.30752e-008              wketa=-5.1334096e-009            pketa=1.6995816e-015 pclm=0.84216358                 lpclm=-1.4301459e-007            wpclm=2.3224719e-008 ppclm=-2.5797631e-014            pdiblc2=0.00041676269              lpdiblc2=7.4813696e-010 wpdiblc2=-4.2585021e-012            ppdiblc2=3.8275416e-017             agidl=1.5939062e-010 lagidl=-3.5063675e-017            wagidl=-5.1907057e-019            pagidl=5.1468269e-024 aigc=0.0067574026               laigc=-2.8816306e-011            waigc=-1.133081e-011 paigc=-6.685944e-018             aigsd=0.0061164928               laigsd=1.7015382e-012 waigsd=-2.7755078e-012            paigsd=2.1708132e-018             tvoff=0.000999914 ltvoff=6.00102e-010               wtvoff=1.19198e-010               ptvoff=-5.64778e-017 kt1=-0.181935                  lkt1=6.9555366e-009             wkt1=3.0749216e-009 pkt1=-6.6792133e-016            kt2=-0.055123402               lkt2=2.7735809e-009 wkt2=8.6205893e-010             pkt2=-7.6550833e-016            ute=-0.93340005 lute=3.6451787e-008             wute=-5.5243993e-010            pute=1.8754954e-015 ua1=2.0432478e-009             lua1=1.2219843e-016             wua1=-4.8094276e-017 pua1=3.0042776e-024             ub1=-2.555872e-018             lub1=1.086231e-025 wub1=1.0191023e-025             pub1=-6.6942565e-032            uc1=3.965463e-010 luc1=2.0740697e-016             wuc1=-2.0663819e-018            puc1=-7.4285611e-024 at=134439.76                  lat=-0.03990453 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=-0.00063111                pat=5.6724167e-009             u0_ff=0.000199677 u0_ss=-0.000199677               u0_sf=0.000110932                u0_fs=-0.000110932 lu0_ff=-1.77314e-10               lu0_ss=1.77314e-10                lu0_sf=-9.85079e-11 lu0_fs=9.85079e-11                wu0_ff=0.0                        wu0_ss=0.0 wu0_sf=4.4e-17                    wu0_fs=-4.4e-17                   pu0_ff=-3.8e-23 pu0_ss=3.8e-23                    pu0_sf=4.5e-23                    pu0_fs=-4.5e-23 ags_ff=-0.0566985                 ags_ss=0.0566985                  ags_sf=-0.023419 ags_fs=0.0624506                  lags_ff=5.03483e-08                lags_ss=-5.03483e-08 lags_sf=2.0796e-08                 lags_fs=-5.54561e-08               wags_ff=6.46363e-09 wags_ss=-6.46363e-09               wags_sf=6.46363e-09                wags_fs=-1.72364e-08 pags_ff=-5.73971e-15               pags_ss=5.73971e-15                pags_sf=-5.73971e-15 pags_fs=1.53059e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.17 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.50834289 lvth0=-3.2205862e-009            wvth0=-8.3319577e-010            pvth0=6.376175e-016 k2=-0.017815342               lk2=-5.9366272e-009            wk2=3.6214873e-009 pk2=-1.6905716e-016            cit=0.0021307482               lcit=-3.7758748e-010 wcit=-1.5756182e-010            pcit=5.2973105e-017             voff=-0.14257764 lvoff=-8.4867585e-009            wvoff=9.8938081e-010             pvoff=3.078569e-016 eta0=0.11407407                 weta0=-3.8844444e-009            etab=-0.063634 wetab=2.139552e-009              u0=0.013358904                lu0=2.0460372e-009 wu0=2.3155368e-010             pu0=-1.5439627e-016            ua=9.4205704e-010 lua=3.2000576e-017             wua=8.1159067e-017             pua=-4.8836358e-023 ub=1.549494e-018              lub=-3.6194153e-025            wub=-1.9649551e-025 pub=9.2946427e-032             uc=-2.4467655e-010            luc=2.833433e-017 wuc=1.2507367e-017             puc=-2.0950195e-024            vsat=133709.63 lvsat=-0.034620818               wvsat=-0.0039310578              pvsat=4.7842993e-009 a0=2.6288929                  la0=-6.9772998e-007            wa0=-8.0575723e-008 pa0=7.5342242e-014             ags=0.66733712                 lags=4.0432691e-007 wags=1.1554439e-008             pags=-1.417376e-014             keta=0.0091908319 lketa=-4.1690699e-009            wketa=-3.7546848e-009            pketa=4.7527397e-016 pclm=1.0408987                  lpclm=-3.1949134e-007            wpclm=-6.5705647e-008 ppclm=5.3172535e-014             pdiblc2=-0.0016571358              lpdiblc2=2.5897588e-009 wpdiblc2=3.6021748e-010             ppdiblc2=-2.8537926e-016            agidl=1.2639695e-010 lagidl=-5.7652939e-018            wagidl=8.1388742e-018             pagidl=-2.541428e-024 aigc=0.0067422413               laigc=-1.5353063e-011            waigc=-1.3882584e-011 paigc=-4.419969e-018             aigsd=0.0061058309               laigsd=1.1169265e-011 waigsd=5.0521378e-012             paigsd=-4.7801361e-018            tvoff=0.00190748 ltvoff=-2.05813e-010              wtvoff=4.42106e-011               ptvoff=1.01113e-017 kt1=-0.16349885                lkt1=-9.4157637e-009            wkt1=3.0012137e-009 pkt1=-6.0246868e-016            kt2=-0.034945058               lkt2=-1.5144788e-008 wkt2=-1.5004234e-009            pkt2=1.3323759e-015             ute=-0.86061467 lute=-2.8181634e-008            wute=7.65624e-009               pute=-5.4138124e-015 ua1=2.5561199e-009             lua1=-3.3323201e-016            wua1=-7.5998936e-017 pua1=2.7783616e-023             ub1=-3.1406344e-018            lub1=6.278921e-025 wub1=1.3272116e-025             pub1=-9.4302669e-032            uc1=5.7962228e-010 luc1=4.48355e-017               wuc1=1.0986692e-017             puc1=-1.9019691e-023 at=179416.78                  lat=-0.079844127 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=-0.0044935129              pat=9.1022305e-009             vsat_ff=576.787 vsat_ss=108.151                    vsat_sf=-2054.81                   vsat_fs=2054.81 lvsat_ff=-0.000512189               lvsat_ss=-9.60359e-05               lvsat_sf=0.00182468 lvsat_fs=-0.00182468                wvsat_ff=0.000378086                wvsat_ss=-0.000567129 wvsat_sf=0.000567129                wvsat_fs=-0.000567129               pvsat_ff=-3.35741e-10 pvsat_ss=5.03611e-10                pvsat_sf=-5.0361e-10                pvsat_fs=5.0361e-10 ags_ff=0.194666                   ags_ss=-0.194666                  lags_ff=-1.72864e-07 lags_ss=1.72864e-07                wags_ff=-7e-15                     wags_ss=7e-15 pags_ff=-3e-20                     pags_ss=3e-20                      at_ff=-8219.26 at_sf=-2054.81                   at_ss=6849.38                    at_fs=2054.81 lat_ff=0.0072987                  lat_sf=0.00182468                 lat_ss=-0.00608225 lat_fs=-0.00182468                wat_ff=0.00226852                 wat_sf=0.000567129 wat_ss=-0.00189043                wat_fs=-0.000567129               pat_ff=-2.01444e-09 pat_sf=-5.0361e-10                pat_ss=1.6787e-09                 pat_fs=5.0361e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.18 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.50191705 lvth0=-6.0351066e-009            wvth0=-6.2636717e-010            pvth0=5.4702657e-016 k2=-0.018703345               lk2=-5.5476821e-009            wk2=2.380136e-009 pk2=3.7465473e-016             cit=0.00082836449              lcit=1.9285657e-010 wcit=9.9404049e-012             pcit=-2.0392869e-017            voff=-0.14677009 lvoff=-6.6504676e-009            wvoff=4.8515081e-010             pvoff=5.2870964e-016 eta0=0.11407407                 weta0=-3.8844444e-009            etab=-0.063634 wetab=2.139552e-009              u0=0.011836643                lu0=2.7127874e-009 wu0=7.2360938e-011             pu0=-8.4669853e-017            ua=1.691777e-009 lua=-2.9637676e-016            wua=-3.8251309e-017            pua=3.465387e-024 ub=4.0510315e-019             lub=1.3930167e-025             wub=2.5061824e-027 pub=5.7836855e-033             uc=-2.3860275e-010            luc=2.5674006e-017 wuc=4.697887e-019              puc=3.1774399e-024             vsat=31708.916 lvsat=0.010055495                wvsat=0.012597109                pvsat=-2.4550377e-009 a0=2.0701804                  la0=-4.5301393e-007            wa0=8.2704536e-008 pa0=3.8254888e-015             ags=-0.96318179                lags=1.1184942e-006 wags=6.1977914e-008             pags=-3.6259243e-014            keta=-0.039003739 lketa=1.6940152e-008             wketa=9.3180701e-009             pketa=-5.2505927e-015 pclm=0.10835728                 lpclm=8.8961782e-008             wpclm=7.884727e-008 ppclm=-1.0141643e-014            pdiblc2=0.0023795821               lpdiblc2=8.2167635e-010 wpdiblc2=-2.0667236e-010            ppdiblc2=-3.7081504e-017            agidl=1.0277033e-010 lagidl=4.5831644e-018             wagidl=1.153426e-018              pagidl=5.181983e-025 aigc=0.0067707018               laigc=-2.7818774e-011            waigc=-2.0951116e-011 paigc=-1.3239521e-018            aigsd=0.0060864958               laigsd=1.9638032e-011 waigsd=-7.6707155e-013            paigsd=-2.2313224e-018            tvoff=0.00131114 ltvoff=5.5382e-011                wtvoff=1.02203e-010               ptvoff=-1.52894e-017 kt1=-0.18716307                lkt1=9.4916413e-010             wkt1=3.4673458e-009 pkt1=-8.0663456e-016            kt2=-0.063820641               lkt2=-2.4972832e-009 wkt2=8.9155303e-010             pkt2=2.8469028e-016             ute=-0.99179584 lute=2.927572e-008              wute=-5.3948957e-009            pute=3.0258508e-016 ua1=1.4720184e-009             lua1=1.4160446e-016             wua1=3.1004928e-017 pua1=-1.9084076e-023            ub1=-2.3406748e-018            lub1=2.775098e-025 wub1=-1.5955735e-025            pub1=3.371532e-032              uc1=4.0881222e-010 luc1=1.1965031e-016             wuc1=-1.8046767e-017            puc1=-6.3030355e-024 at=32404.627                  lat=-0.015452804 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=0.026073587                pat=-4.2861591e-009            vsat_ff=279.196 vsat_ss=-4825.25                   vsat_sf=884.137                    vsat_fs=-2111.11 lvsat_ff=-0.000381848               lvsat_ss=0.0020648                  lvsat_sf=0.00053741 lvsat_fs=-3.4e-10                   wvsat_ff=-0.000388447               wvsat_ss=0.000921309 wvsat_sf=-0.000244022               wvsat_fs=0.000582667                pvsat_ff=3e-17 pvsat_ss=-1.48326e-10               pvsat_sf=-1.48326e-10               pvsat_fs=-3e-17 ags_ff=-0.374359                  ags_ss=0.374359                   lags_ff=7.63697e-08 lags_ss=-7.63697e-08               wags_ff=-3.2e-14                   wags_ss=3.2e-14 pags_ff=2e-21                      pags_ss=-2e-21                     at_ff=15806.3 at_sf=3951.57                    at_ss=-13171.9                   at_fs=-3951.57 lat_ff=-0.00322448                lat_sf=-0.00080612                lat_ss=0.00268707 lat_fs=0.00080612                 wat_ff=-0.00436253                wat_sf=-0.00109063 wat_ss=0.00363544                 wat_fs=0.00109063                 pat_ff=8.89956e-10 pat_sf=2.22489e-10                pat_ss=-7.4163e-10                pat_fs=-2.22489e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.19 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.5294396 lvth0=-4.2050692e-010            wvth0=2.6543525e-009             pvth0=-1.2224024e-016 k2=-0.030933017               lk2=-3.0528291e-009            wk2=5.0490939e-009 pk2=-1.6981269e-016            cit=0.00087199602              lcit=1.8395574e-010 wcit=-1.1024237e-010            pcit=4.1244168e-018             voff=-0.16011228 lvoff=-3.9286603e-009            wvoff=2.2143223e-009             pvoff=1.7595866e-016 eta0=0.11407407                 weta0=-3.8844444e-009            etab=-0.063633981 wetab=2.1395499e-009             u0=0.022689312                lu0=4.9884297e-010 wu0=-3.3668787e-010            pu0=-1.2238949e-018            ua=7.3647291e-10 lua=-1.0149473e-16             wua=-6.1998607e-17             pua=8.3098358e-24 ub=6.2891491e-019             lub=9.364407e-026              wub=1.1133633e-025 pub=-1.6417665e-032            uc=-2.8251199e-010            luc=3.463149e-017 wuc=3.5116081e-017             puc=-3.8904036e-024            vsat=73297.377 lvsat=0.0015714486               wvsat=0.0010244566               pvsat=-9.4216624e-011 a0=1.751538                   la0=-3.8801086e-007            wa0=2.6634621e-007 pa0=-3.3637413e-014            ags=5.0247319                  lags=-1.030402e-007 wags=-6.7193768e-008            pags=-9.9082194e-015            keta=0.20932143 lketa=-3.3718183e-008            wketa=-2.5382643e-008            pketa=1.8283528e-015 pclm=0.62400353                 lpclm=-1.6230053e-008            wpclm=4.4763598e-008 ppclm=-3.188574e-015             pdiblc2=0.008952381                lpdiblc2=-5.191746e-010 wpdiblc2=-7.4914286e-010            ppdiblc2=7.3582476e-017             agidl=1.4559112e-010 lagidl=-4.1522768e-018            wagidl=-2.1214042e-018            pagidl=1.1862637e-024 aigc=0.0067324762               laigc=-2.0020741e-011            waigc=-2.4456967e-011 paigc=-6.0875837e-019            aigsd=0.0061573383               laigsd=5.1861636e-012 waigsd=-9.1275933e-012            paigsd=-5.2577598e-019            tvoff=0.00240687 ltvoff=-1.68146e-010              wtvoff=-9.03865e-011              ptvoff=2.39989e-017 kt1=-0.14222729                lkt1=-8.2177358e-009            wkt1=-3.7290061e-009 pkt1=6.6142123e-016             kt2=-0.080776074               lkt2=9.6162522e-010 wkt2=3.1067581e-009             pkt2=-1.6721156e-016            ute=-0.83787355 lute=-2.1244269e-009            wute=-1.6458698e-008            pute=2.5596008e-015 ua1=1.9690123e-009             lua1=4.021771e-017              wua1=-2.5056743e-017 pua1=-7.6474954e-024            ub1=-4.8286771e-019            lub1=-1.0148285e-025 wub1=-6.8305973e-026            pub1=1.5100039e-032             uc1=1.3426777e-009 luc1=-7.0858256e-017            wuc1=-7.5717174e-017            puc1=5.4617275e-024 at=-95798.807                 lat=0.010700696 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=0.010249638                pat=-1.0580735e-009            letab=-3.8297312e-015 petab=4.3658936e-022             vsat_ff=-2761.9                    vsat_ss=6465.59 vsat_sf=5696.65                    vsat_fs=-4724.87                   lvsat_ff=0.000238539 lvsat_ss=-0.00023854                lvsat_sf=-0.000444339               lvsat_fs=0.000533206 wvsat_ff=-0.000749141               wvsat_ss=0.000554925                wvsat_sf=-0.00157228 wvsat_fs=0.00130406                 pvsat_ff=7.35825e-11                pvsat_ss=-7.35825e-11 pvsat_sf=1.22637e-10                pvsat_fs=-1.47165e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_12_mac.20 pmos ( level=54                         lmin=6.299e-08                  lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.57182308 lvth0=2.8854047e-009             wvth0=4.8746913e-009             pvth0=-2.9542667e-016 k2=2.6267395e-005             lk2=-5.4676533e-009            wk2=1.1797548e-009 pk2=1.3199576e-016             cit=0.0029137966               lcit=2.4695296e-011 wcit=-6.7358797e-011            pcit=7.7949801e-019             voff=-0.21863585 lvoff=6.3617834e-010             wvoff=9.7089668e-009             pvoff=-4.0862361e-016 eta0=0.11407407                 weta0=-3.8844444e-009            etab=-0.12987778 wetab=8.953826e-009              u0=0.03455908                 lu0=-4.269989e-010 wu0=-4.8618679e-010            pu0=1.0437021e-017             ua=-6.6853642e-10 lua=8.0959968e-18              wua=5.1786721e-17              pua=-5.6541982e-25 ub=1.9538229e-018             lub=-9.6987501e-027            wub=-9.1084845e-026 pub=-6.2881302e-034            uc=3.3197119e-010             luc=-1.3298198e-017 wuc=-3.0536049e-017            puc=1.2304625e-024             vsat=110614.18 lvsat=-0.0013392614              wvsat=-0.0025817146              pvsat=1.8706473e-010 a0=7.3276617                  la0=-8.2294852e-007            wa0=-8.6583387e-007 pa0=5.4672633e-014             ags=3.7037037                  lags=0 wags=-1.9422222e-007            pags=0                          keta=-0.26773663 lketa=3.4923457e-009             wketa=-3.1291358e-008            pketa=2.2892326e-015 pclm=0.62497662                 lpclm=-1.6305954e-008            wpclm=-2.774688e-008 ppclm=2.4672433e-015             pdiblc2=0.0036255144               lpdiblc2=-1.0367901e-010 wpdiblc2=-1.7264198e-010            ppdiblc2=2.8615407e-017             agidl=1.8493862e-011 lagidl=5.7613093e-018             wagidl=5.3115365e-018             pagidl=6.0649429e-025 aigc=0.0066048263               laigc=-1.0064052e-011            waigc=-3.0871037e-011 paigc=-1.0846098e-019            aigsd=0.006264601                laigsd=-3.1803197e-012 waigsd=2.3349046e-011             paigsd=-3.0589539e-018            tvoff=-0.00165421 ltvoff=1.48618e-010               wtvoff=4.60977e-010               ptvoff=-1.90075e-017 kt1=-0.27330254                lkt1=2.0061339e-009             wkt1=8.2852843e-009 pkt1=-2.7569343e-016            kt2=-0.08880695                lkt2=1.5880336e-009 wkt2=-1.7339967e-010            pkt2=8.8640749e-017             ute=-1.1437534 lute=2.1734201e-008             wute=3.8081073e-008             pute=-1.6945014e-015 ua1=2.5144218e-009             lua1=-2.3242351e-018            wua1=-1.5801737e-016 pua1=2.7234336e-024             ub1=-1.2584257e-018            lub1=-4.0989331e-026 wub1=8.7264151e-026             pub1=2.9655691e-033             uc1=3.0386608e-010 luc1=1.0169052e-017             wuc1=9.2281949e-018             puc1=-1.1640113e-024 at=62658.728                  lat=-0.0016589913 jtsswgs='1e-009*(1+1200*0.06*iboffp_flag_12)'                              jtsswgd='1e-009*(1+1200*0.06*iboffp_flag_12)' wat=-0.0070251822              pat=2.8936242e-010             letab=5.1670123e-009 petab=-5.315131e-016             vsat_ff=-5576.92                   vsat_ss=16272.5 vsat_fs=6096.51                    vsat_mc=2573.03                    lvsat_ff=0.000458111 lvsat_ss=-0.00100348                lvsat_fs=-0.000310861               lvsat_mc=-0.000200696 wvsat_ff=0.00129419                 wvsat_ss=-0.00185507                wvsat_fs=-0.00168264 wvsat_mc=-0.000293325               pvsat_ff=-8.57976e-11               pvsat_ss=1.14397e-10 pvsat_fs=8.57976e-11                pvsat_mc=2.28794e-11 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_18_mac.global nmos ( modelid=9                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=0                          igbmod=0 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_18'              permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=3.36e-009                  toxm=3.36e-009                  dtox=2.83e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=1e-008 xw=0                          dlc=1.17e-008                  dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.31 k3=-5.1                       k3b=0.25                       w0=0 dvt0=0.0103                     dvt1=0.02                       dvt2=-0.09 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.4                       voffl=-5e-009 dvtp0=1.5e-006                   dvtp1=0                          lpe0=8e-008 lpeb=5e-009                     xj=6.7e-008                   ngate=4.8e+020 ndep=1e+017                     nsd=1e+020                     phin=0.15 cdsc=0                          cdscb=0                          cdscd=0 ud=0                          nfactor=0.7                        a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=0.45 delta=0.01                       pscbe1=9.264e+008                 pscbe2=1e-020 fprout=750                        pdits=0                          pditsd=0 pditsl=0                          rsh=18.0                       rdsw=150 prwg=0                          prwb=0                          wr=1 alpha0=0                          alpha1=0.06                       beta0=8.83 bgidl=1.1e+009                   cgidl=5                          egidl=0.8 aigbacc=0.01238                    bigbacc=0.006109                   cigbacc=0.2809 nigbacc=4.05                       aigbinv=0.35                       bigbinv=0.03 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1 aigc=0.009898                   bigc=0.001383                   cigc=1.515e-005 aigsd=0.0086                     bigsd=0.0004353                  cigsd=3.925e-020 nigc=1                          poxedge=1                          pigcd=1.672 ntox=1                          cgso=4.5e-011                   cgdo=4.5e-011 cgbo=0                          cgdl=7.9e-011                   cgsl=7.9e-011 clc=0                          cle=0.6                        cf='8.09e-011+5.742e-11*ccoflag_18' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=5                          noff=3                          voffcv=-0.085 kt1l=0                          kt2=-0.03                      prt=0 fnoimod=1                          tnoimod=1                          em=2.53e+009 ef=0.94                       noia=0                          noib=0 noic=0                          lintnoi=-3.80e-008                 jss=2.69e-07 jsd=2.69e-07                   jsws=7.06e-14                   jswd=7.06e-14 jswgs=7.06e-14                   jswgd=7.06e-14                   njs=1.09 njd=1.09                       ijthsfwd=0.01                       ijthdfwd=0.01 ijthsrev=0.01                       ijthdrev=0.01                       bvs=7.9 bvd=7.9                        xjbvs=1                          xjbvd=1 jtsswgs=2e-009                     jtsswgd=2e-009                     njtsswg=15 xtsswgs=0.5                        xtsswgd=0.5                        tnjtsswg=1 vtsswgs=1                          vtsswgd=1                          pbs=0.715 pbd=0.715                      cjs=0.001472                   cjd=0.001472 mjs=0.336                      mjd=0.336                      pbsws=0.457 pbswd=0.457                      cjsws=1.086e-010                 cjswd=1.086e-010 mjsws=0.015                      mjswd=0.015                      pbswgs=0.923 pbswgd=0.923                      cjswgs=2.016e-010                 cjswgd=2.016e-010 mjswgs=0.552                      mjswgd=0.552                      tpb=0.00137 tcj=0.00079                    tpbsw=0.00230                    tcjsw=0.00020 tpbswg=0.00114                    tcjswg=0.00073                    xtis=3 xtid=3                          dmcg=6.7e-008                   dmci=6.7e-008 dmdg=0                          dmcgt=0                          dwj=0 xgw=0                          xgl=2.64e-009                  rshg=16.42 gbmin=1e-012                     rbpb=50                         rbpd=50 rbps=50                         rbdb=50                         rbsb=50 ngcon=1                          xrcrg1=12                         xrcrg2=1 pk2we=0                          lk2we=0                          wk2we=0 k2we=0                          pku0we=-1e-16                     wku0we=0 lku0we=0                          ku0we=-0.004                     pkvth0we=-1e-17 wkvth0we=0                          lkvth0we=0                          kvth0we=0.0085 wec=-2800                      web=-150                       scref=1e-6 wpemod=1                          rnoia=0                          rnoib=0 tnoia=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.5 sigma_factor='sigma_factor_18' ccoflag='ccoflag_18' rcoflag='rcoflag_18' rgflag='rgflag_18' mismatchflag='mismatchflag_mos_18' globalflag='globalflag_mos_18' totalflag='totalflag_mos_18' global_factor='global_factor_18' local_factor='local_factor_18' sigma_factor_flicker='sigma_factor_flicker_18' noiseflag='noiseflagn_18' noiseflag_mc='noiseflagn_18_mc' delvto=0 mulu0=1 dlc_fmt=2 par1_io='par1_io' par2_io='par2_io' par3_io='par3_io' par4_io='par4_io' par5_io='par5_io' par6_io='par6_io' par7_io='par7_io' par8_io='par8_io' par9_io='par9_io' par10_io='par10_io' par11_io='par11_io' par12_io='par12_io' par13_io='par13_io' par14_io='par14_io' par15_io='par15_io' par16_io='par16_io' par17_io='par17_io' par18_io='par18_io' par19_io='par19_io' par20_io='par20_io' w1_io='2.0857*0.40825' w2_io='0.67082*-0.40825' w3_io='0.54772*0.26807' w4_io='0.54772*-0.6902' w5_io='0.54772*-0.32981' w6_io='0.54772*0.098267' tox_c='toxn_18'                  dxl_c='dxln_18'                  dxw_c='dxwn_18' ddlc_c='ddlcn_18'                 cgo_c='cgon_18'                  cgl_c='cgln_18' cj_c='cjn_18'                   cjsw_c='cjswn_18'                 cjswg_c='cjswgn_18' cf_c='cfn_18'                   dvth_c='dvthn_18'                 dwvth_c='dwvthn_18' dlvth_c='dlvthn_18'                dpvth_c='dpvthn_18'                du0_c='du0n_18' dwu0_c='dwu0n_18'                 dlu0_c='dlu0n_18'                 dpu0_c='dpu0n_18' dk2_c='dk2n_18'                  dwk2_c='dwk2n_18'                 dlk2_c='dlk2n_18' dpk2_c='dpk2n_18'                 dags_c='dagsn_18'                 dwags_c='dwagsn_18' dpdiblc2_c='dpdiblc2n_18'             dlpdiblc2_c='dlpdiblc2n_18'            dvsat_c='dvsatn_18' dwvsat_c='dwvsatn_18'               duc_c='ducn_18'                  dluc_c='dlucn_18' dwuc_c='dwucn_18'                 dpuc_c='dpucn_18'                 dketa_c='dketan_18' dlketa_c='dlketan_18'               dwketa_c='dwketan_18'               dpketa_c='dpketan_18' monte_flag_c='monte_flagn_18'          c1f_c='c1fn_18'                  c2f_c='c2fn_18' c3f_c='c3fn_18' global_mc='global_mc_flag_18' tox_g='toxn_18_ms_global'        dxl_g='dxln_18_ms_global'        dxw_g='dxwn_18_ms_global' cgo_g='cgon_18_ms_global'        cgl_g='cgln_18_ms_global'        cj_g='cjn_18_ms_global' cjsw_g='cjswn_18_ms_global'       cjswg_g='cjswgn_18_ms_global'      cf_g='cfn_18_ms_global' dvth_g='dvthn_18_ms_global'       dwvth_g='dwvthn_18_ms_global'      dlvth_g='dlvthn_18_ms_global' dpvth_g='dpvthn_18_ms_global'      du0_g='du0n_18_ms_global'        dwu0_g='dwu0n_18_ms_global' dlu0_g='dlu0n_18_ms_global'       dpu0_g='dpu0n_18_ms_global'       dk2_g='dk2n_18_ms_global' dwk2_g='dwk2n_18_ms_global'       dlk2_g='dlk2n_18_ms_global'       dpk2_g='dpk2n_18_ms_global' dags_g='dagsn_18_ms_global'       dwags_g='dwagsn_18_ms_global'      dvsat_g='dvsatn_18_ms_global' dwvsat_g='dwvsatn_18_ms_global'     dluc_g='dlucn_18_ms_global'       dlketa_g='dlketan_18_ms_global' monte_flag_g='monte_flagn_18_ms_global' weight1=2.2047059 weight2=-1.8575882 weight3=-0.90158824 weight4=-0.58823529 weight5=-0.40471765 tox_1=-2.3955414e-011 tox_2=-8.9373236e-012 tox_3=-1.6291481e-012 tox_4=9.4219297e-011 tox_5=5.1583358e-013 dxl_1=-1.4376247e-009 dxl_2=-5.3637536e-010 dxl_3=-9.7773875e-011 dxl_4=-5.6546372e-009 dxl_5=3.0957612e-011 dxl_max=-2.2e-008 dxw_1=7.0729697e-010 dxw_2=-2.6725306e-009 dxw_3=-7.8365641e-010 dxw_4=4.2997794e-025 dxw_5=-1.1643341e-008 dxw_max=-1.2e-008 cgo_1=3.7272e-013 cgo_2=-2.2768e-013 cgo_3=-6.1739e-014 cgo_4=-2.8927e-029 cgo_5=7.9899e-014 cgl_1=6.5432e-013 cgl_2=-3.9971e-013 cgl_3=-1.0839e-013 cgl_4=-2.848e-029 cgl_5=1.4027e-013 cj_1=-1.2192e-005 cj_2=7.4477e-006 cj_3=2.0195e-006 cj_4=7.2531e-022 cj_5=-2.6136e-006 cjsw_1=-8.9949e-013 cjsw_2=5.4947e-013 cjsw_3=1.49e-013 cjsw_4=3.1935e-029 cjsw_5=-1.9282e-013 cjswg_1=-1.6698e-012 cjswg_2=1.02e-012 cjswg_3=2.7659e-013 cjswg_4=5.9716e-029 cjswg_5=-3.5795e-013 cf_1=6.7006e-013 cf_2=-4.0932e-013 cf_3=-1.1099e-013 cf_4=-1.9574e-029 cf_5=1.4364e-013 dvth_1=-0.0017428 dvth_2=0.008148 dvth_3=0.0018262 dvth_4=-3.0783e-019 dvth_5=-0.0020616 dwvth_1=-6.5967e-010 dwvth_2=7.2666e-010 dwvth_3=6.096e-011 dwvth_4=-9.2199e-027 dwvth_5=-2.0574e-010 dlvth_1=-2.158761e-010 dlvth_2=3.345166e-010 dlvth_3=8.974691e-011 dlvth_4=3.283335e-028 dlvth_5=-9.395166e-011 dpvth_1=4.6949e-017 dpvth_2=4.1044e-017 dpvth_3=2.2304e-017 dpvth_4=-1.1223e-032 dpvth_5=-6.5162e-018 du0_1=0.00015496 du0_2=0.00028363 du0_3=5.1554e-005 du0_4=-2.3503e-021 du0_5=-5.9431e-005 dwu0_1=7.763e-011 dwu0_2=9.4157e-011 dwu0_3=-6.7442e-012 dwu0_4=-6.9556e-027 dwu0_5=-1.6664e-011 dlu0_1=2.1018e-011 dlu0_2=2.2904e-011 dlu0_3=-1.9334e-012 dlu0_4=-2.8615e-027 dlu0_5=-3.5708e-012 dpu0_1=1.1718e-017 dpu0_2=5.39912e-018 dpu0_3=-8.6297e-019 dpu0_4=3.7638e-034 dpu0_5=-9.3827e-019 dk2_1=0.0004774 dk2_2=0.00094815 dk2_3=0.00018641 dk2_4=-7.4278e-020 dk2_5=-0.00019284 dwk2_1=-7.3502e-012 dwk2_2=3.9212e-012 dwk2_3=1.1925e-011 dwk2_4=4.8506e-028 dwk2_5=-2.2095e-012 dlk2_1=3.3952e-011 dlk2_2=7.7131e-011 dlk2_3=1.2768e-011 dlk2_4=-1.1238e-026 dlk2_5=-1.6938e-011 dpk2_1=-4.101e-018 dpk2_2=2.8935e-018 dpk2_3=-6.6306e-018 dpk2_4=-8.8094e-034 dpk2_5=-4.4646e-019 dags_1=0.0021372 dags_2=0.0029623 dags_3=-0.0027687 dags_4=5.229e-019 dags_5=-0.00038734 dwags_1=-2.9389e-009 dwags_2=-1.1743e-009 dwags_3=-6.8702e-010 dwags_4=6.9762e-025 dwags_5=7.139e-011 dvsat_1=51.986 dvsat_2=-15.831 dvsat_3=-308.43 dvsat_4=-1.1821e-014 dvsat_5=28.89 dwvsat_1=7.4621e-005 dwvsat_2=3.73695e-005 dwvsat_3=-4.2311e-005 dwvsat_4=1.1036e-020 dwvsat_5=-1.6368e-005 dluc_1=-1.7928e-019 dluc_2=1.3227e-019 dluc_3=-3.9862e-019 dluc_4=3.9001e-035 dluc_5=-1.3081e-020 dlketa_1=8.9641e-011 dlketa_2=-6.6135e-011 dlketa_3=1.9931e-010 dlketa_4=-1.4829e-026 dlketa_5=6.5405e-012 monte_flag_1=-0.179775 monte_flag_2=-0.0670738 monte_flag_3=-0.0122266 monte_flag_4=-0.707113 monte_flag_5=0.00387125 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.9998 b_4=-0.0009597                 c_4=-0.00141                   d_4=-0.001335 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.0035                     mis_a_2=-0.0405                    mis_a_3=0.0339 mis_b_1=0.001                      mis_b_2=0                          mis_b_3=0 mis_c_1=0.5                        mis_c_2=0                          mis_c_3=0 mis_d_1=0.00087                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.0061                     mis_e_2=-0.076                     mis_e_3=0.0329 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=0                          xl0=1e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0                       bidirectionflag=1 designflag=1 cf0=8.09e-011                  cco=5.742e-11 noimod=6                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718                      tnoiamax=9593223.1145 tnoiac1=123552.3055                tnoiac2=9231959.0635               rnoiamax=0.61424 rnoiac1=0.0085845                  rnoiac2=0.58914 saref0=0.468e-6            sbref0=0.468e-6 samax=10e-6               sbmax=10e-6 samin=0.135e-6            sbmin=0.135e-6 rllodflag=0                   lreflod=1e-6                llodref=1 lod_clamp=-1e90 wlod0=0 ku00=0e-9                lku00=0e-15               wku00=0e-15 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=0 kvth00=-0e-10            lkvth00=-0e-16              wkvth00=-0e-16 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                 lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=3e-9                lku000=1e-15               wku000=1e-15       		pku000=0 llodku000=1                   wlodku000=1 kvth000=-2.5e-10              lkvth000=-3e-16            wkvth000=-6e-16     		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0.2                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=-1e-7               lku01=-1.5e-14            wku01=2e-14 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0.2 kvth01=2e-8                lkvth01=3e-22               wkvth01=3e-15 pkvth01=4.5e-29             llodvth1=2                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=-0.15               lodk21=1 wlod2=0 ku02=0                   lku02=0                   wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0 kvth02=0                   lkvth02=0                   wkvth02=0 pkvth02=0                   llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0                   lku03=0                   wku03=0 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0 kvth03=0                   lkvth03=0                   wkvth03=0 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=0                   lku003=0                   wku003=0         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=4.68e-7             sa_b1=1.35e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.98e-7             spamax=1.6e-6              spamin=1.98e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=0.01                wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl=0.8e-10             ldplkvth0=1.36                pkvth0dpl=0.0e-19 ku0dpl=0.0                 wku0dpl=0e-8                wdplku0=1 lku0dpl=3.2e-6              ldplku0=0.8                 pku0dpl=0.0e-11 keta0dpl=0.5                 wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0.5                 wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx=-0.0                wku0dpx=0e-9                wdpxku0=1 lku0dpx=0.0e-8              ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=0.00                wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps=0.0                 wku0dps=-0.0e-9             wdpsku0=1 lku0dps=0.0e-16             ldpsku0=1.0                 pku0dps=0.0e-23 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=-0.00               wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa=0.0e-9              ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa=0.00                wku0dpa=0e-7                wdpaku0=1 lku0dpa=0.0e-11             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=-0.0                wka0dpa=0                   wdpaka0=1 lka0dpa=-0.0e-7             ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=1.0                 wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.31e-7             spbmax='1.6e-6+1.6e-6+0.135e-6'    spbmin='1.98e-7+1.98e-7+0.135e-6' pse_mode=1 kvth0dp2=0.004               wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0.7e-8              ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.000               wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=0.35e-5             ldp2ku0=0.7                 pku0dp2=0 keta0dp2=0.1                 wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0.8                 wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=1.0                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=10e-6               enxmax=10e-6		 enxmin=0.18e-6 kvth0enx='0.010*3'           wkvth0enx='0.7e-8*2'          wenxkvth0=1 lkvth0enx='4e-5*0'            lenxkvth0=1.0                 pkvth0enx=-3.3e-16 ku0enx='-0.60-0.2'         wku0enx='-0.8e-7*1'         wenxku0=1 lku0enx='0.2e-7'            lenxku0=1                   pku0enx=-3.7e-15 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx='0.0-1'             wka0enx=0                   wenxka0=1 lka0enx='1.0e-7*0'          lenxka0=1.0                 pka0enx='1.0e-14*0' kvsatenx='0.65*1'            wenx=0                   ku0enx0='0.10' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.045e-6 kvth0eny='0.01'              wkvth0eny='3.5e-8*1'          wenykvth0=1 lkvth0eny='1e-7*0'            lenykvth0=1.0                 pkvth0eny=0 ku0eny='(-0.5)*1'          wku0eny='(-0.2e-7)*1'       wenyku0=1 ku0eny0='0.41+0.01'         wku0eny0='-1e-7*2'           weny0ku0=1 lku0eny='(1.2e-11)*1'       lenyku0='1.5'               pku0eny='5.0e-19*0' keta0eny=0.00                wketa0eny=0                   wenyketa0=1 ka0eny='-0.50*1'           wka0eny='-2e-7*0'           wenyka0=1 lka0eny='-6.0e-8*0'         lenyka0=1.0                 pka0eny='(1.0e-14)*0' kvsateny='-0.6+0.4'          weny=1e-6 kvth0eny1=0.000              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=0 ku0eny1='(0.15)*0'         wku0eny1=0.0e-8             weny1ku0=1 lku0eny1='0.0e-5'           leny1ku0=1.0                pku0eny1=-0.0e-14 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1.0                pka0eny1=0 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=2e-5	         ringxmax=9.027e-6		 ringxmin=4.770e-07 kvth0rx=-0.1                wkvth0rx=-1.0e-8             wrxkvth0=1.0 lkvth0rx=0.0e-9              lrxkvth0=1.0                 pkvth0rx=0.0e-16 ku0rx=1.00                wku0rx=1.0e-8              wrxku0=1.0 lku0rx='1.0e-7'            lrxku0=1.0                 pku0rx=0.0e-15 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.0                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=12e-6               ringymax=9.027e-6		 ringymin=0.477e-6 kvth0ry='-0.005'            wkvth0ry='-1e-8*5'           wrykvth0=1.0 lkvth0ry=0.0e-8              lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry=0.1                 wku0ry='1.0e-7*0.3'        wryku0=1.0 lku0ry='1e-5*1'            lryku0=1                   pku0ry=-0.0e-16 keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry=0.0                 wry=1e-6 kvth0ry0=-0.00               ku0ry0=0.01 sfxref=1.89e-7           sfxmax=3e-6               minwodx=0.53e-6 sfxmin=0.189e-6 lrefodx=5e-8              lodxref=1                 wodx=1e-6 kvth0odxa=-0.200            lkvth0odxa=1.0e-13           lodxakvth0=2.0 wkvth0odxa=1.0e-11           wodxakvth0=2.0               pkvth0odxa=0.0e-16 ku0odxa=-0.30             lku0odxa=3.0e-13           lodxaku0=2.0 wku0odxa=5.0e-11           wodxaku0=2.0               pku0odxa=-0.0e-26 keta0odx=0.10              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0005           lkvth0odx1b=0.0e-7            lodx1bkvth0=0.5 wkvth0odx1b=-0.0e-15          wodx1bkvth0=2.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.001            lku0odx1b=0.0e-7            lodx1bku0=0.5 wku0odx1b=-0.5e-14          wodx1bku0=2.0               pku0odx1b=0.0e-16 sfyref=8.1e-7 sfymin=0.15e-6 sfymax=3e-6              minwody=0e-7              wody=1e-6 kvth0odya=-0.000            lkvth0odya=1.0e-13           lodyakvth0=2.0 wkvth0odya=0.0e-6            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=-2.00             lku0odya=2.0e-13           lodyaku0=2.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=0.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.00             lkvth0odyb=-3.0e-9           lodybkvth0=1.0 wkvth0odyb=-7.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=0.10              lku0odyb=0.0e-9            lodybku0=0.8 wku0odyb=-0.0e-5           wodybku0=1.0               pku0odyb=0.0e-13 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_18_mac.1 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-006                     wmax=0.00090001                 vth0=0.43516 k2=0.014574632                cit=0.0015                     voff=-0.17146719 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.5470274e-009            ub=2.510615e-018              uc=1.01528e-010 vsat=100000                     a0=1.8                        ags=0.77816907 keta=-0.060714323               pclm=0.2365                     pdiblc2=0.001 agidl=4.7909339e-010             tvoff=0.001815                   kt1=-0.198016 ute=-1                         ua1=2.2203714e-009             ub1=-2.08e-018 uc1=-3.5e-011                  at=120000                     lvth0=0 lk2=0                          luc=0                          lketa=0 lpdiblc2=0                          lu0=0                          wvth0=0 wk2=0                          wuc=0                          wags=0 wketa=0                          pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18_mac.2 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-006                     wmax=0.00090001                 vth0=0.43583426 k2=0.01610097                 cit=0.0015550505               voff=-0.17176577 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.5479495e-009            ub=2.5120759e-018             uc=1.0290646e-010 vsat=100275.25                  a0=1.8421412                  ags=0.71539931 keta=-0.058904163               pclm=0.17959154                 pdiblc2=0.0009583364 agidl=5.1730707e-010             tvoff=0.00183644                 kt1=-0.19457754 ute=-1                         ua1=2.2881347e-009             ub1=-2.1212879e-018 uc1=-3.6238636e-011            at=121126.33                  lvth0=-6.0750761e-009 lk2=-1.3752307e-008            lcit=-4.9600505e-010            lvoff=2.6902347e-009 lua=8.3079606e-018             lub=-1.3162734e-026            luc=-1.2419966e-017 lvsat=-0.0024800252              la0=-3.7969187e-007            lags=5.6555552e-007 lketa=-1.6309534e-008            lpclm=5.1274522e-007             lpdiblc2=3.7538902e-010 lagidl=-3.4430524e-016            ltvoff=-1.93194e-010              lkt1=-3.0980476e-008 lua1=-6.1054678e-016            lub1=3.7200379e-025             luc1=1.1160114e-017 lat=-0.010148263               lu0=0                          wvth0=0 wk2=0                          wuc=0                          wags=0 wketa=0                          pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18_mac.3 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-006                     wmax=0.00090001                 vth0=0.42963686 k2=0.0074962214               cit=0.0011                     voff=-0.16750235 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.4981584e-009            ub=2.5566613e-018             uc=9.36624e-011 vsat=98000                      a0=1.7875156                  ags=0.80265184 keta=-0.064214382               pclm=0.65                       pdiblc2=0.00031105711 agidl=2.9517105e-010             tvoff=0.0017434                  kt1=-0.2102 ute=-1                         ua1=1.641984e-009              ub1=-1.5524444e-018 uc1=-1.32e-011                 at=194043.2                   lvth0=6.8009024e-010 lk2=-4.3731311e-009            lvoff=-1.9568951e-009            lua=-4.5964306e-017 lub=-6.1760853e-026            luc=-2.343936e-018             la0=-3.2014996e-007 lags=4.7045026e-007             lketa=-1.0521396e-008            lpdiblc2=1.0809234e-009 lagidl=-1.0217698e-016            ltvoff=-9.17732e-011              lkt1=-1.3952e-008 lua1=9.375744e-017              lub1=-2.4803556e-025            luc1=-1.3952e-017 lat=-0.089627648               lu0=0                          wvth0=0 wk2=0                          wuc=0                          wags=0 wketa=0                          pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18_mac.4 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-006                     wmax=0.00090001                 vth0=0.43995888 k2=0.0052985221               cit=0.000944                   voff=-0.1757704 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.6427414e-009            ub=2.6595534e-018             uc=9.2652e-011 vsat=98503.496                  a0=2.6980475                  ags=0.66058977 keta=-0.1215324                 pclm=0.728                      pdiblc2=-0.00018914922 agidl=1.2975302e-010             tvoff=0.00173603                 kt1=-0.21162952 ute=-0.688                     ua1=2.7247733e-009             ub1=-2.4704e-018 uc1=-3.5e-011                  at=97009.2                    lvth0=-5.9260032e-009 lk2=-2.9666036e-009            lcit=9.984e-011                 lvoff=3.334656e-009 lua=4.656883e-017              lub=-1.2761174e-025            luc=-1.69728e-018 lvsat=-0.00032223759             la0=-9.0289038e-007            lags=5.6136999e-007 lketa=2.6162136e-008             lpclm=-4.992e-008                lpdiblc2=1.4010555e-009 lagidl=3.6905546e-018             ltvoff=-8.70605e-011              lkt1=-1.3037107e-008 lua1=-5.992277e-016             lub1=3.39456e-025               lat=-0.027525888 lute=-1.9968e-007               lu0=0                          wvth0=0 wk2=0                          wuc=0                          wags=0 wketa=0                          pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18_mac.5 nmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=9e-006                     wmax=0.00090001                 vth0=0.42400175 k2=-0.0041934273              cit=0.00084489796              voff=-0.17859039 eta0=0.18                       etab=-0.035                     u0=0.019857143 ua=-1.6888162e-009            ub=2.2035268e-018             uc=8.137551e-011 vsat=99853.575                  a0=1.5873206                  ags=2.277551 keta=-0.056962347               pclm=0.68877551                 pdiblc2=0.0042338257 agidl=6.1972392e-011             tvoff=0.00101524                 kt1=-0.25633722 ute=-1.2                       ua1=1.5469318e-009             ub1=-1.777551e-018 uc1=-4.9795918e-011            at=25175.832                  lvth0=2.9727943e-010 lk2=7.3525667e-010             lcit=1.384898e-010              lvoff=4.4344523e-009 lua=6.4537988e-017             lub=5.0238616e-026             luc=2.700551e-018 lvsat=-0.00084876841             la0=-4.6970691e-007            lags=-6.9244898e-008 lketa=9.7981531e-010             lpclm=-3.4622449e-008            lpdiblc2=-3.2390473e-010 lagidl=3.0125e-017                ltvoff=1.94047e-010               lkt1=4.3988975e-009 lua1=-1.3986951e-016            lub1=6.9244898e-026             luc1=5.7704082e-018 lat=0.00048912553              lu0=1.6157143e-009             wvth0=0 wk2=0                          wuc=0                          wags=0 wketa=0                          pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18_mac.6 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-007                     wmax=9e-006                     vth0=0.43536861 k2=0.014923896                cit=0.0015362917               voff=-0.17107143 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.5469007e-009            ub=2.5162389e-018             uc=1.0250889e-010 vsat=100000                     a0=1.7667745                  ags=0.77929598 keta=-0.061386044               pclm=0.23777778                 pdiblc2=0.00099777778 agidl=4.8625058e-010             tvoff=0.00184031                 kt1=-0.19767822 ute=-1                         ua1=2.229546e-009              ub1=-2.0944444e-018 uc1=-3.625e-011                at=120000                     lvth0=0 lk2=0                          luc=0                          lketa=0 lpdiblc2=0                          lu0=0                          wvth0=-1.8775e-009 wk2=-3.1433799e-009            wcit=-3.26625e-010              wvoff=-3.56181e-009 weta0=-1.6e-007                  wetab=-5e-009                    wua=-1.1406e-018 wub=-5.0615e-026               wuc=-8.828e-018                wa0=2.9902927e-007 wags=-1.0142204e-008            wketa=6.04549e-009               wpclm=-1.15e-008 wpdiblc2=2e-011                     wagidl=-6.4414719e-017            wtvoff=-2.278e-010 wkt1=-3.04e-009                 wua1=-8.257142e-017             wub1=1.3e-025 wuc1=1.125e-017                 pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.7 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-007                     wmax=9e-006                     vth0=0.43590596 k2=0.01649581                 cit=0.001597866                voff=-0.17133744 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.5483953e-009            ub=2.5176355e-018             uc=1.0396895e-010 vsat=100275.25                  a0=1.8060001                  ags=0.71664671 keta=-0.059691733               pclm=0.1787514                  pdiblc2=0.00095758632 agidl=5.253547e-010              tvoff=0.00186195                 kt1=-0.19437984 ute=-1                         ua1=2.2996729e-009             ub1=-2.1387907e-018 uc1=-3.7721836e-011            at=121089.39                  lvth0=-4.8414984e-009 lk2=-1.4162942e-008            lcit=-5.5478509e-010            lvoff=2.3967598e-009 lua=1.3466952e-017             lub=-1.2583373e-026            luc=-1.3155156e-017 lvsat=-0.0024800252              la0=-3.5342229e-007            lags=5.6446997e-007 lketa=-1.526574e-008             lpclm=5.3182764e-007             lpdiblc2=3.6212502e-010 lagidl=-3.5232809e-016            ltvoff=-1.94944e-010              lkt1=-2.9718418e-008 lua1=-6.318435e-016             lub1=3.9955962e-025             luc1=1.3261246e-017 lat=-0.0098153888              lu0=0                          wvth0=-6.4529147e-010 wk2=-3.5535595e-009            wcit=-3.853398e-010             wvoff=-3.8549592e-009 weta0=-1.6e-007                  wetab=-5e-009                    wua=4.0126654e-018 wub=-5.0036282e-026            wuc=-9.5623737e-018            wa0=3.2526969e-007 wags=-1.1226547e-008            wketa=7.0881252e-009             wpclm=7.5612374e-009 wpdiblc2=6.7507197e-012             wagidl=-7.242866e-017             wtvoff=-2.29548e-010 wkt1=-1.7793434e-009            wua1=-1.0384451e-016            wub1=1.5752525e-025 wuc1=1.3348801e-017             pvth0=-1.1102199e-014            pk2=3.6957182e-015 pcit=5.2902039e-016             pvoff=2.641274e-015              pua=-4.6430921e-023 pub=-5.2142531e-033            puc=6.6167074e-024             pa0=-2.3642619e-013 pags=9.769928e-015              pketa=-9.3941432e-015            ppclm=-1.7174175e-013 ppdiblc2=1.1937602e-016             pagidl=7.220561e-023              ptvoff=1.57482e-017 pkt1=-1.1358516e-014            pua1=1.9167051e-022             pub1=-2.4800252e-031 puc1=-1.8910193e-023            wat=0.00033250505              pat=-2.9958705e-009 wvsat=0                          wu0=0                          pu0=0 pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.8 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-007                     wmax=9e-006                     vth0=0.43133578 k2=0.0069306501               cit=0.0010730864               voff=-0.16930915 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.485957e-009             ub=2.5603284e-018             uc=9.2971407e-011 vsat=98000                      a0=1.7524593                  ags=0.78149618 keta=-0.061446508               pclm=0.71407407                 pdiblc2=0.00013786191 agidl=2.9400029e-010             tvoff=0.0017208                  kt1=-0.20691654 ute=-1                         ua1=1.6023032e-009             ub1=-1.495679e-018 uc1=-1.0385185e-011            at=192442.77                  lvth0=1.3999437e-010 lk2=-3.7369182e-009            lcit=1.7224691e-011             lvoff=1.8592332e-010 lua=-5.4590802e-017            lub=-5.9118586e-026            luc=-1.1678341e-018 la0=-2.9506285e-007            lags=4.9378405e-007             lketa=-1.3353035e-008 lpclm=-5.1674074e-008            lpdiblc2=1.2556246e-009             lagidl=-1.0015178e-016 ltvoff=-4.10981e-011              lkt1=-1.6053412e-008            lua1=1.282895e-016 lub1=-3.014321e-025             luc1=-1.6535704e-017            lat=-0.08759057 lu0=0                          wvth0=-1.5290302e-008            wk2=5.090142e-009 wcit=2.4222222e-010             wvoff=1.6261224e-008             weta0=-1.6e-007 wetab=-5e-009                    wua=-1.0981246e-016            wub=-3.3003111e-026 wuc=6.2189333e-018             wa0=3.1550616e-007             wags=1.9040097e-007 wketa=-2.4910859e-008            wpclm=-5.7666667e-007            wpdiblc2=1.5587568e-009 wagidl=1.0536865e-017             wtvoff=2.03318e-010               wkt1=-2.9551111e-008 wua1=3.5712711e-016             wub1=-5.1088889e-025            wuc1=-2.5333333e-017 pvth0=4.8608628e-015             pk2=-5.7259164e-015            pcit=-1.5502222e-016 pvoff=-1.9285366e-014            pua=7.7638462e-023             pub=-2.3780409e-032 puc=-1.0584917e-023            pa0=-2.2578395e-013            pags=-2.1000406e-013 pketa=2.548475e-014              ppclm=4.6506667e-013             ppdiblc2=-1.5723107e-015 pagidl=-1.8226812e-023            ptvoff=-4.56075e-016              pkt1=1.8912711e-014 pua1=-3.1078855e-022            pub1=4.8056889e-031             puc1=2.3253333e-023 wat=0.014403911                pat=-1.8333703e-008            wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.9 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-007                     wmax=9e-006                     vth0=0.4417723 k2=0.0054507845               cit=0.00096133333              voff=-0.17468974 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.6498193e-009            ub=2.6739037e-018             uc=9.3575283e-011 vsat=98559.44                   a0=2.787875                   ags=0.63581794 keta=-0.12567426                pclm=0.70266667                 pdiblc2=-3.6296727e-006 agidl=1.3617223e-010             tvoff=0.00183725                 kt1=-0.20953947 ute=-0.65333333                ua1=2.7936121e-009             ub1=-2.5144e-018 uc1=-3.3795556e-011            at=99058.349                  lvth0=-6.5393762e-009 lk2=-2.7898043e-009            lcit=8.8746667e-011             lvoff=3.629499e-009 lua=5.0281044e-017             lub=-1.3180683e-025            luc=-1.5543147e-018 lvsat=-0.00035804177             la0=-9.5772887e-007            lags=5.8701812e-007 lketa=2.7752725e-008             lpclm=-4.4373333e-008            lpdiblc2=1.3461792e-009 lagidl=8.5817738e-019             ltvoff=-1.15626e-010              lkt1=-1.4374741e-008 lua1=-6.3414818e-016            lub1=3.5054933e-025             luc1=-1.5530667e-018 lat=-0.027824544               lute=-2.2186667e-007            lu0=0 wvth0=-1.6320762e-008            wk2=-1.3703621e-009            wcit=-1.56e-010 wvoff=-9.7259296e-009            weta0=-1.6e-007                  wetab=-5e-009 wua=6.3700638e-017             wub=-1.2915335e-025            wuc=-8.30955e-018 wa0=-8.0844748e-007            wags=2.2294652e-007             wketa=3.7276713e-008 wpclm=2.28e-007                  wpdiblc2=-1.6696759e-009            wagidl=-5.7772834e-017 wtvoff=-9.11e-010                 wkt1=-1.881048e-008             wua1=-6.1954928e-016 wub1=3.96e-025                  wuc1=-1.084e-017                pvth0=5.5203573e-015 pk2=-1.5911938e-015            pcit=9.984e-017                 pvoff=-2.6535875e-015 pua=-3.3409919e-023            pub=3.7755744e-032             puc=-1.286688e-024 pa0=4.9354638e-013             pags=-2.3083321e-013            pketa=-1.4315296e-014 ppclm=-4.992e-014                ppdiblc2=4.938863e-016              pagidl=2.5491395e-023 ptvoff=2.57088e-016               pkt1=1.2038707e-014             pua1=3.1428434e-022 pub1=-9.984e-032                puc1=1.39776e-023               wat=-0.018442343 pat=2.6878995e-009             wvsat=-0.00050349624             pvsat=3.2223759e-010 wute=-3.12e-007                 pute=1.9968e-013                wu0=0 pu0=0                          u0_mc=3.46667e-05                lu0_mc=-2.21867e-11 wu0_mc=-3.12e-10                  pu0_mc=1.9968e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.10 nmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=9e-007                     wmax=9e-006                     vth0=0.42462821 k2=-0.0036779275              cit=0.00083837687              voff=-0.17771724 eta0=0.19777778                 etab=-0.034444444               u0=0.019857143 ua=-1.6811312e-009            ub=2.188862e-018              uc=8.0798373e-011 vsat=99665.553                  a0=1.4576238                  ags=2.3362286 keta=-0.056688151               pclm=0.68752834                 pdiblc2=0.0048541029 agidl=5.5747575e-011             tvoff=0.00101335                 kt1=-0.25720893 ute=-1.1959184                 ua1=1.5820317e-009             ub1=-1.8023129e-018 uc1=-5.1455782e-011            at=26962.815                  lvth0=1.4681734e-010 lk2=7.7039341e-010             lcit=1.3669969e-010             lvoff=4.8102244e-009 lua=6.2492687e-017             lub=5.735946e-026              luc=3.4286804e-018 lvsat=-0.00078942563             la0=-4.3893092e-007            lags=-7.6142036e-008 lketa=8.4814293e-010             lpclm=-3.8469388e-008            lpdiblc2=-5.4833644e-010 lagidl=3.2223791e-017             ltvoff=2.05697e-010               lkt1=4.2163475e-009 lua1=-1.6163183e-016            lub1=7.2835374e-026             luc1=5.3344218e-018 lat=0.00029271504              lute=-1.0258503e-008            lu0=1.6157143e-009 wvth0=-5.638202e-009             wk2=-4.6394984e-009            wcit=5.8689796e-011 wvoff=-7.8583354e-009            weta0=-1.6e-007                  wetab=-5e-009 wua=-6.9165066e-017            wub=1.3198342e-025             wuc=5.1942347e-018 wa0=1.1672712e-006             wags=-5.2809826e-007            wketa=-2.4677684e-009 wpclm=1.122449e-008              wpdiblc2=-5.5824941e-009            wagidl=5.6023357e-017 wtvoff=1.70418e-011               wkt1=7.8453061e-009             wua1=-3.1589958e-016 wub1=2.2285714e-025             wuc1=1.4938776e-017             pvth0=1.3541588e-015 pk2=-3.1623067e-016            pcit=1.611098e-017              pvoff=-3.3819492e-015 pua=1.8407706e-023             pub=-6.4087596e-032            puc=-6.553164e-024 pa0=-2.7698391e-013            pags=6.2074247e-014             pketa=1.1850514e-015 ppclm=3.4622449e-014             ppdiblc2=2.0198854e-015             pagidl=-1.8889119e-023 ptvoff=-1.04848e-016              pkt1=1.6429506e-015             pua1=1.9586096e-022 pub1=-3.2314286e-032            puc1=3.9238775e-024             wat=-0.016082843 pat=1.7676944e-009             wvsat=0.0016922029               pvsat=-5.3408509e-010 wute=-3.6734694e-008            pute=9.2326531e-014             wu0=0 pu0=0                          u0_mc=-2.22223e-05               vsat_mc=-131.519 lvsat_mc=5.12925e-05                lu0_mc=-1.7e-18                   wvsat_mc=0.00118367 pvsat_mc=-4.61633e-10               wu0_mc=2e-10                      pu0_mc=-3.5e-23 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.11 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=5.4e-007                   wmax=9e-007                     vth0=0.44265375 k2=0.015628011                cit=0.0002773125               voff=-0.19156542 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.477435e-009             ub=2.4e-018                   uc=9.945e-011 vsat=100000                     a0=2.0975732                  ags=0.75891614 keta=-0.060655368               pclm=0.2625                     pdiblc2=0.001025238 agidl=3.6634794e-010             tvoff=0.000855116                kt1=-0.19975742 ute=-1                         ua1=1.845236e-009              ub1=-1.425e-018 uc1=-2.375e-012                at=120000                     lvth0=0 lk2=0                          luc=0                          lketa=0 lpdiblc2=0                          lu0=0                          wvth0=-8.434125e-009 wk2=-3.7770834e-009            wcit=8.0645625e-010             wvoff=1.4882778e-008 weta0=1.755e-007                 wetab=7.7274e-009                wua=-6.3659722e-017 wub=5.4e-026                   wuc=-6.075e-018                wa0=1.3104855e-009 wags=8.1996584e-009             wketa=5.3878817e-009             wpclm=-3.375e-008 wpdiblc2=-4.7142e-012               wagidl=4.3497655e-017             wtvoff=6.58876e-010 wkt1=-1.168722e-009             wua1=2.6330762e-016             wub1=-4.725e-025 wuc1=-1.92375e-017              pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.12 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=0.44529752 k2=0.016742369                cit=0.00012968253              voff=-0.1948109 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.4690192e-009            ub=2.3947771e-018             uc=9.9373205e-011 vsat=100275.25                  a0=2.1756294                  ags=0.67913341 keta=-0.055751144               pclm=0.26077967                 pdiblc2=0.00078132821 agidl=3.8013043e-010             tvoff=0.000736711                kt1=-0.19432055 ute=-1                         ua1=1.8143026e-009             ub1=-1.304577e-018 uc1=4.5235164e-012             at=119088.91                  lvth0=-2.3820333e-008 lk2=-1.0040366e-008            lcit=1.330146e-009              lvoff=2.9241755e-008 lua=-7.5825805e-017            lub=4.7058479e-026             luc=6.9192705e-019 lvsat=-0.0024800252              la0=-7.0328661e-007            lags=7.1884237e-007 lketa=-4.4187057e-008            lpclm=1.5500158e-008             lpdiblc2=2.1976273e-009 lagidl=-1.2418024e-016            ltvoff=1.06683e-009               lkt1=-4.8986178e-008 lua1=2.7871022e-016             lub1=-1.085011e-024             luc1=-6.2155633e-017 lat=0.0082088836               lu0=0                          wvth0=-9.0976935e-009 wk2=-3.775463e-009             wcit=9.3602536e-010             wvoff=1.7271149e-008 weta0=1.755e-007                 wetab=7.7274e-009                wua=-6.7425822e-017 wub=6.0536284e-026             wuc=-5.4262023e-018            wa0=-7.3966958e-009 wags=2.2535422e-008             wketa=3.5415951e-009             wpclm=-6.6264205e-008 wpdiblc2=1.6538302e-010             wagidl=5.8273177e-017             wtvoff=7.83165e-010 wkt1=-1.8327029e-009            wua1=3.3298884e-016             wub1=-5.9326705e-025 wuc1=-2.4672017e-017            pvth0=5.9787519e-015             pk2=-1.4599933e-017 pcit=-1.1674176e-015            pvoff=-2.1519221e-014            pua=3.393256e-023 pub=-5.889192e-032             puc=-5.8456675e-024            pa0=7.8451704e-014 pags=-1.2916523e-013            pketa=1.6635042e-014             ppclm=2.9295298e-013 ppdiblc2=-1.532576e-015             pagidl=-1.3312746e-022            ptvoff=-1.11984e-015 pkt1=5.9824682e-015             pua1=-6.2782784e-022            pub1=1.0881111e-030 puc1=4.8964999e-023             wat=0.0021329318               pat=-1.9217716e-008 wvsat=0                          wu0=0                          pu0=0 pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.13 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=0.41687939 k2=0.015027069                cit=0.0014922222               voff=-0.14124298 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.6691786e-009            ub=2.5914789e-018             uc=1.1317493e-010 vsat=98000                      a0=2.6758876                  ags=1.3561141 keta=-0.13521583                pclm=-0.57833333                pdiblc2=0.0071245349 agidl=4.6390646e-010             tvoff=0.00266137                 kt1=-0.25058004 ute=-1                         ua1=2.3680978e-009             ub1=-2.8333333e-018 uc1=-8.45e-011                 at=268625.78                  lvth0=7.1554227e-009 lk2=-8.1706889e-009            lcit=-1.5502222e-010            lvoff=-2.9147278e-008 lua=1.4234791e-016             lub=-1.6734649e-025            luc=-1.4351957e-017 la0=-1.2485681e-006            lags=-1.9066563e-008            lketa=4.2429448e-008 lpclm=9.3013333e-007             lpdiblc2=-4.716468e-009             lagidl=-2.154961e-016 ltvoff=-1.03105e-009              lkt1=1.2336668e-008             lua1=-3.2492658e-016 lub1=5.8133333e-025             luc1=3.488e-017                 lat=-0.1547863 lu0=0                          wvth0=-2.2795517e-009            wk2=-2.1966346e-009 wcit=-1.35e-010                 wvoff=-8.9983344e-009            weta0=1.755e-007 wetab=7.7274e-009                wua=5.5086963e-017             wub=-6.10386e-026 wuc=-1.196424e-017             wa0=-5.1557932e-007            wags=-3.2675515e-007 wketa=4.1481528e-008             wpclm=5.865e-007                 wpdiblc2=-4.7292488e-009 wagidl=-1.4237869e-016            wtvoff=-6.43191e-010              wkt1=9.74604e-009 wua1=-3.32088e-016              wub1=6.93e-025                  wuc1=4.137e-017 pvth0=-1.4530227e-015            pk2=-1.7355228e-015            pcit=-1.8994406e-030 pvoff=7.1145155e-015             pua=-9.9606377e-023            pub=7.3624704e-032 puc=1.2807936e-024             pa0=6.3237077e-013             pags=2.5156149e-013 pketa=-2.4719484e-014            ppclm=-4.1856e-013               ppdiblc2=3.8025727e-015 pagidl=8.5583078e-023             ptvoff=4.34884e-016               pkt1=-6.6383616e-015 pua1=9.710592e-023              pub1=-3.1392e-031               puc1=-2.30208e-023 wat=-0.0541608                 pat=4.2142452e-008             wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.14 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.42823758 k2=0.0074162525               cit=0.000704                   voff=-0.18830252 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.3845577e-009            ub=2.3768e-018                uc=8.6293031e-011 vsat=98000                      a0=0.335                      ags=0.82358353 keta=-0.076892699               pclm=1.148                      pdiblc2=-0.0053070628 agidl=3.7786914e-011             tvoff=0.000364301                kt1=-0.23801824 ute=-1                         ua1=2.6341272e-009             ub1=-2.627e-018 uc1=-5.652e-011                at=48359.117                  lvth0=-1.138176e-010 lk2=-3.2997666e-009            lcit=3.4944e-010                lvoff=9.7083018e-010 lua=-3.9809478e-017            lub=-2.9952e-026               luc=2.85246e-018 la0=2.496e-007                 lags=3.2175299e-007             lketa=5.1026455e-009 lpclm=-1.7472e-007               lpdiblc2=3.2397545e-009             lagidl=5.7220404e-017 ltvoff=4.39071e-010               lkt1=4.2971136e-009             lua1=-4.9518543e-016 lub1=4.4928e-025                luc1=1.69728e-017               lat=-0.013815635 lu0=0                          wvth0=-4.139516e-009             wk2=-3.1392832e-009 wcit=7.56e-011                  wvoff=2.5255733e-009             weta0=1.755e-007 wetab=7.7274e-009                wua=-1.750348e-016             wub=1.3824e-025 wuc=-1.7555231e-018            wa0=1.39914e-006               wags=5.3957483e-008 wketa=-6.6266894e-009            wpclm=-1.728e-007                wpdiblc2=3.1034139e-009 wagidl=3.0773946e-017             wtvoff=4.14658e-010               wkt1=6.820416e-009 wua1=-4.7601292e-016            wub1=4.9734e-025                wuc1=9.612e-018 pvth0=-2.6264549e-016            pk2=-1.1322277e-015            pcit=-1.34784e-016 pvoff=-2.6078548e-016            pua=4.7671551e-023             pub=-5.39136e-032 puc=-5.2527852e-024            pa0=-5.930496e-013             pags=7.9054051e-015 pketa=6.0697748e-015             ppclm=6.7392e-014                ppdiblc2=-1.2103314e-015 pagidl=-2.5234608e-023            ptvoff=-2.42139e-016              pkt1=-4.7659622e-015 pua1=1.8921787e-022             pub1=-1.886976e-031             puc1=-2.69568e-024 wat=0.027186966                pat=-9.9201184e-009            wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0                          u0_mc=-0.000312                  lu0_mc=1.9968e-10 wu0_mc=0.0                        pu0_mc=0.0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.15 nmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.4278394 k2=0.0016137502               cit=0.00087529592              voff=-0.1893543 eta0=-0.175                     etab=-0.048586                  u0=0.019857143 ua=-1.7426736e-009            ub=2.4242857e-018             uc=1.1704793e-010 vsat=106164.86                  a0=3.8942246                  ags=0.99673701 keta=-0.075270054               pclm=0.54020408                 pdiblc2=-0.0080268894 agidl=1.9167852e-010             tvoff=0.00132648                 kt1=-0.24353592 ute=-1.5918367                 ua1=4.6462701e-010             ub1=-1.3122449e-018 uc1=-6.0938775e-011            at=7534.9734                  lvth0=4.1472154e-011 lk2=-1.0367907e-009            lcit=2.8263459e-010             lvoff=1.3810247e-009 lua=9.9855737e-017             lub=-4.8471429e-026            luc=-9.1419495e-018 lvsat=-0.003184294               la0=-1.1384976e-006            lags=2.5422313e-007 lketa=4.4698141e-009             lpclm=6.2320408e-008             lpdiblc2=4.3004868e-009 lagidl=-2.7973237e-018            ltvoff=6.38207e-011               lkt1=6.4490082e-009 lua1=3.5091965e-016             lub1=-6.347449e-026             luc1=1.8696122e-017 lat=0.0021057812               lute=2.3081633e-007             lu0=1.6157143e-009 wvth0=-8.5282722e-009            wk2=-9.4020082e-009            wcit=2.5462653e-011 wvoff=2.6150196e-009             weta0=1.755e-007                 wetab=7.7274e-009 wua=-1.3776875e-017            wub=-7.9897959e-026            wuc=-2.7430364e-017 wa0=-1.0256695e-006            wags=6.7744418e-007             wketa=1.4255945e-008 wpclm=1.4381633e-007             wpdiblc2=6.0103989e-009             wagidl=-6.6314496e-017 wtvoff=-2.64778e-010              wkt1=-4.4604e-009               wua1=6.8976465e-016 wub1=-2.1820408e-025            wuc1=2.3473469e-017             pvth0=1.4489694e-015 pk2=1.310235e-015              pcit=-1.1523044e-016            pvoff=-2.9566952e-016 pua=-1.5219039e-023            pub=3.1160204e-032             puc=4.7604028e-024 pa0=3.5262611e-013             pags=-2.3525441e-013            pketa=-2.0744527e-015 ppclm=-5.6088367e-014            ppdiblc2=-2.3440556e-015            pagidl=1.2629884e-023 ptvoff=2.28404e-017               pkt1=-3.66444e-016              pua1=-2.6543538e-022 pub1=9.0364592e-032             puc1=-8.1016531e-024            wat=0.0014022142 pat=1.359349e-010              wvsat=-0.0041571703              pvsat=1.6212964e-009 wute=3.1959184e-007             pute=-1.2464082e-013            wu0=0 pu0=0                          u0_mc=2.2449e-05                 vsat_mc=1627.55 lvsat_mc=-0.000634743               lu0_mc=6.92451e-11                wvsat_mc=-0.000399491 pvsat_mc=1.55801e-10                wu0_mc=1.59796e-10                pu0_mc=-6.23204e-17 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.16 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.42910039 k2=0.016243241                cit=0.00135265                 voff=-0.1681236 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.6175468e-009            ub=2.62e-018                  uc=1.0786e-010 vsat=100000                     a0=2.3                        ags=0.87190207 keta=-0.07279409                pclm=0.2                        pdiblc2=0.001133524 agidl=6.4044621e-010             tvoff=0.00209897                 kt1=-0.20486516 ute=-1                         ua1=2.764928e-009              ub1=-2.9e-018 uc1=-5.8e-011                  at=120000                     lvth0=0 lk2=0                          luc=0                          lketa=0 lpdiblc2=0                          lu0=0                          wvth0=-1.1153117e-009 wk2=-4.1093078e-009            wcit=2.25774e-010               wvoff=2.2241952e-009 weta0=-8.64e-008                 wetab=1.001808e-008              wua=1.200069e-017 wub=-6.48e-026                 wuc=-1.06164e-017              wa0=-1.08e-007 wags=-5.2812744e-008            wketa=1.1942791e-008             wpdiblc2=-6.318864e-011 wagidl=-1.0451541e-016            wtvoff=-1.28045e-011              wkt1=1.5894576e-009 wua1=-2.3332609e-016            wub1=3.24e-025                  wuc1=1.08e-017 pvth0=0                          pk2=0                          puc=0 pketa=0                          wvsat=0                          wu0=0 pu0=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.17 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.43046267 k2=0.016946903                cit=0.001359896                voff=-0.16659847 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.6215494e-009            ub=2.6441204e-018             uc=1.0860848e-010 vsat=100275.25                  a0=2.3756944                  ags=0.85336935 keta=-0.073629861               pclm=0.16240051                 pdiblc2=0.0011381378 agidl=7.2765024e-010             tvoff=0.00224871                 kt1=-0.19934563 ute=-1                         ua1=2.9306917e-009             ub1=-3.1050631e-018 uc1=-6.4479444e-011            at=124475.61                  lvth0=-1.2274131e-008 lk2=-6.3399888e-009            lcit=-6.5286665e-011            lvoff=-1.3741403e-008 lua=3.6062828e-017             lub=-2.1732461e-025            luc=-6.7438087e-018 lvsat=-0.0024800252              la0=-6.8200694e-007            lags=1.6697981e-007 lketa=7.5302965e-009             lpclm=3.3877145e-007             lpdiblc2=-4.1570183e-011 lagidl=-7.8570829e-016            ltvoff=-1.34919e-009              lkt1=-4.9731004e-008 lua1=-1.4935308e-015            lub1=1.8476188e-024             luc1=5.8379794e-017 lat=-0.040325211               lu0=0                          wvth0=-1.0868769e-009 wk2=-3.8859112e-009            wcit=2.7171007e-010             wvoff=2.0364389e-009 weta0=-8.64e-008                 wetab=1.001808e-008              wua=1.4940457e-017 wub=-7.4109096e-026            wuc=-1.0413251e-017            wa0=-1.1543182e-007 wags=-7.1551984e-008            wketa=1.3196102e-008             wpclm=-1.3139454e-008 wpdiblc2=-2.7294147e-011            wagidl=-1.2938752e-016            wtvoff=-3.33155e-011 wkt1=8.8083671e-010             wua1=-2.6986131e-016            wub1=3.7899545e-025 wuc1=1.2589582e-017             pvth0=-2.5619692e-016            pk2=-2.0128038e-015 pcit=-4.1388397e-016            pvoff=1.6916839e-015             pua=-2.6487302e-023 pub=8.387495e-032              puc=-1.8303702e-024            pa0=6.6960682e-014 pags=1.6884055e-013             pketa=-1.1292329e-014            ppclm=1.1838649e-013 ppdiblc2=-3.2340938e-016            pagidl=2.2409769e-022             ptvoff=1.84804e-016 pkt1=6.3846742e-015             pua1=3.291823e-022              pub1=-4.9550905e-031 puc1=-1.6124132e-023            wat=-0.00077588182             pat=6.9906952e-009 wvsat=0                          wu0=0                          pu0=0 pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.18 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.40825089 k2=0.026188636                cit=0.0023170222               voff=-0.14985865 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.5635028e-009            ub=2.3803702e-018             uc=1.2319627e-010 vsat=98000                      a0=1.9633333                  ags=0.22111143 keta=-0.057600561               pclm=0.50619556                 pdiblc2=-0.00018 agidl=-2.0011244e-010            tvoff=0.00155439                 kt1=-0.26821861 ute=-1                         ua1=1.5935893e-009             ub1=-1.0686667e-018 uc1=5.4688666e-012             at=121763.2                   lvth0=1.1936711e-008 lk2=-1.6413478e-008            lcit=-1.1085542e-009            lvoff=-3.1987806e-008 lua=-2.7207919e-017            lub=7.0163058e-026             luc=-2.2644499e-017 la0=-2.3253333e-007            lags=8.5614093e-007             lketa=-9.9416399e-009 lpclm=-3.5965156e-008            lpdiblc2=1.3952e-009                lagidl=2.2555302e-016 ltvoff=-5.92375e-010              lkt1=2.5340552e-008             lua1=-3.6089173e-017 lub1=-3.7205333e-025            luc1=-1.7863865e-017            lat=-0.037368688 lu0=0                          wvth0=2.37984e-009               wk2=-8.2238811e-009 wcit=-5.8039199e-010            wvoff=-4.3458699e-009            weta0=-8.64e-008 wetab=1.001808e-008              wua=-1.9779576e-018            wub=5.296008e-026 wuc=-1.7375762e-017            wa0=-1.308e-007                wags=2.8614629e-007 wketa=-4.307161e-010             wpclm=8.544e-010                 wpdiblc2=-7.848e-010 wagidl=2.1619151e-016             wtvoff=-4.54198e-011              wkt1=1.9270867e-008 wua1=8.614656e-017              wub1=-2.5992e-025               wuc1=-7.2131879e-018 pvth0=-4.0349184e-015            pk2=2.7155834e-015             pcit=5.1490727e-016 pvoff=8.6484006e-015             pua=-8.04623e-024              pub=-5.4630451e-032 puc=5.7587661e-024             pa0=8.3712e-014                pags=-2.2105056e-013 pketa=3.5609032e-015             ppclm=1.0313318e-013             ppdiblc2=5.02272e-016 pagidl=-1.5258345e-022            ptvoff=1.97998e-016               pkt1=-1.3660459e-014 pua1=-5.8866278e-023            pub1=2.009088e-031              puc1=5.4608869e-024 wat=0.025144992                pat=-2.1263057e-008            wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0                          u0_mc=0.000284444                lu0_mc=-3.10044e-10 wu0_mc=-1.536e-10                 pu0_mc=1.67424e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.19 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.42382441 k2=0.011945321                cit=-3.7094974e-005            voff=-0.20219733 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.6241451e-009            ub=2.6928e-018                uc=1.0987428e-010 vsat=98000                      a0=2.146                      ags=2.0811878 keta=-0.09597384                pclm=0.4032                     pdiblc2=-0.00268 agidl=3.2981508e-010             tvoff=0.000731214                kt1=-0.21719232 ute=-1                         ua1=2.0848255e-009             ub1=-2.43e-018 uc1=-6.993516e-011             at=142692.69                  lvth0=1.9696595e-009 lk2=-7.2977563e-009            lcit=3.9808079e-010             lvoff=1.5089478e-009 lua=1.1603155e-017             lub=-1.29792e-025              luc=-1.4118427e-017 la0=-3.4944e-007               lags=-3.3430793e-007            lketa=1.4617258e-008 lpclm=2.9952e-008                lpdiblc2=2.9952e-009                lagidl=-1.1360058e-016 ltvoff=-6.5545e-011               lkt1=-7.3162752e-009            lua1=-3.5048033e-016 lub1=4.992e-025                 luc1=3.0394712e-017             lat=-0.050763563 lu0=0                          wvth0=-1.7564026e-009            wk2=-5.5849801e-009 wcit=4.7579129e-010             wvoff=1.002877e-008              weta0=-8.64e-008 wetab=1.001808e-008              wua=-4.5657581e-017            wub=-3.24e-026 wuc=-1.4489399e-017            wa0=4.212e-007                 wags=-6.2514881e-007 wketa=3.6771267e-009             wpclm=2.29392e-007               wpdiblc2=1.6848e-009 wagidl=-1.2692126e-016            wtvoff=2.16525e-010               wkt1=-4.4255808e-009 wua1=-1.7938999e-016            wub1=3.9096e-025                wuc1=1.6856186e-017 pvth0=-1.3877231e-015            pk2=1.0266867e-015             pcit=-1.6105003e-016 pvoff=-5.51369e-016              pua=1.9908729e-023             pub=-1.7913775e-045 puc=3.9114937e-024             pa0=-2.69568e-013              pags=3.621783e-013 pketa=9.3188385e-016             ppclm=-4.313088e-014             ppdiblc2=-1.078272e-015 pagidl=6.7008726e-023             ptvoff=3.03534e-017               pkt1=1.5052677e-015 pua1=1.1107711e-022             pub1=-2.156544e-031             puc1=-9.9435127e-024 wat=-0.023753164               pat=1.0031763e-008             wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0                          u0_mc=-0.000824                  lu0_mc=3.9936e-10 wu0_mc=2.7648e-10                 pu0_mc=-1.07827e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.20 nmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.42673106 k2=-0.0093237196              cit=0.001092301                voff=-0.20711602 eta0=0.31                       etab=-0.052828                  u0=0.019857143 ua=-1.641151e-009             ub=2.1469388e-018             uc=6.8745074e-011 vsat=98200.608                  a0=1.8721589                  ags=1.8300216 keta=-0.073219292               pclm=0.66938775                 pdiblc2=0.010515236 agidl=-5.3456526e-011            tvoff=0.000157831                kt1=-0.24776033 ute=-0.52653061                ua1=2.5336766e-009             ub1=-1.7122449e-018 uc1=2.6086531e-011             at=2788.9622                  lvth0=8.3606567e-010 lk2=9.971694e-010              lcit=-4.2383648e-011            lvoff=3.4272386e-009 lua=1.8235438e-017             lub=8.3093878e-026             luc=1.9219643e-018 lvsat=-7.823704e-005             la0=-2.4264198e-007            lags=-2.3635314e-007 lketa=5.7429849e-009             lpclm=-7.3861224e-008            lpdiblc2=-2.1509422e-009 lagidl=3.5875339e-017             ltvoff=1.58075e-010               lkt1=4.6052474e-009 lua1=-5.2553226e-016            lub1=2.1927551e-025             luc1=-7.0537469e-018 lat=0.0037988918               lute=-1.8465306e-007            lu0=1.6157143e-009 wvth0=-7.9297669e-009            wk2=-3.4957746e-009            wcit=-9.1720102e-011 wvoff=1.220635e-008              weta0=-8.64e-008                 wetab=1.001808e-008 wua=-6.8599102e-017            wub=6.9869388e-026             wuc=-1.3468234e-018 wa0=6.6245972e-008             wags=2.2747047e-007             wketa=1.3148534e-008 wpclm=7.4057143e-008             wpdiblc2=-4.002349e-009             wagidl=6.605843e-017 wtvoff=3.66294e-010               wkt1=-2.1792196e-009            wua1=-4.2752214e-016 wub1=-2.2040816e-027            wuc1=-2.3520196e-017            pvth0=1.0198889e-015 pk2=2.1189658e-016             pcit=6.0279415e-017             pvoff=-1.400625e-015 pua=2.8855922e-023             pub=-3.9885061e-032            puc=-1.2141106e-024 pa0=-1.3113593e-013            pags=2.9656782e-014             pketa=-2.7619649e-015 ppclm=1.7449714e-014             ppdiblc2=1.1397161e-015             pagidl=-8.2533537e-024 ptvoff=-2.80566e-017              pkt1=6.2918684e-016             pua1=2.0784865e-022 pub1=-6.2320408e-032            puc1=5.8032764e-024             wat=0.0039650602 pat=-7.783448e-010             wvsat=0.0001435239               pvsat=-5.5974321e-011 wute=-2.5567347e-007            pute=9.9712653e-014             wu0=0 pu0=0                          u0_mc=0.000318367                vsat_mc=2071.43 lvsat_mc=-0.000807854               lu0_mc=-4.61635e-11               wvsat_mc=-0.000639184 pvsat_mc=2.49281e-10                wu0_mc=-2.7e-16                   pu0_mc=-2.7e-23 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.21 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.39330752 k2=0.0076464838               cit=0.002299                   voff=-0.15436512 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-1.865698e-009             ub=2.4e-018                   uc=5.4471019e-011 vsat=100000                     a0=1.2                        ags=0.572 keta=-0.03187431                pclm=0.30304                    pdiblc2=0.000838 agidl=-5.41322e-013              tvoff=0.0023061                  kt1=-0.21177 ute=-1                         ua1=1.7432e-009                ub1=-1.68e-018 uc1=-1.2e-011                  at=120000                     lvth0=0 lk2=0                          luc=0                          lketa=0 lpdiblc2=0                          lu0=0                          wvth0=1.1770122e-008 wk2=-1.0144751e-009            wcit=-1.14912e-010              wvoff=-2.7288576e-009 weta0=1.152e-007                 wetab=1.4688e-008                wua=1.013351e-016 wub=1.44e-026                  wuc=8.6036332e-018             wa0=2.88e-007 wags=5.5152e-008                wketa=-2.7883292e-009            wpclm=-3.70944e-008 wpdiblc2=4.32e-011                  wagidl=1.262401e-016              wtvoff=-8.7372e-011 wkt1=4.0752e-009                wua1=1.34496e-016               wub1=-1.152e-025 wuc1=-5.76e-018                 pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=2.88e-009                  pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.22 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.39272144 k2=0.0096380468               cit=0.0024777765               voff=-0.14973871 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-1.8291497e-009            ub=2.3637836e-018             uc=5.488193e-011 vsat=100275.25                  a0=1.0098155                  ags=0.54445742 keta=-0.0310503                 pclm=0.16693313                 pdiblc2=0.0013662096 agidl=-3.6673871e-011            tvoff=0.00259595                 kt1=-0.20323417 ute=-1                         ua1=1.8738701e-009             ub1=-1.842399e-018 uc1=-1.6789394e-011            at=116404.45                  lvth0=5.280569e-009 lk2=-1.7943983e-008            lcit=-1.6107764e-009            lvoff=-4.1683917e-008 lua=-3.2929969e-016            lub=3.2630932e-025             luc=-3.7023136e-018 lvsat=-0.0024800252              la0=1.7135619e-006             lags=2.4815862e-007 lketa=-7.4243277e-009            lpclm=1.2263229e-006             lpdiblc2=-4.7591685e-009 lagidl=3.2555427e-016             ltvoff=-2.61158e-009              lkt1=-7.6907865e-008 lua1=-1.1773374e-015            lub1=1.4632149e-024             luc1=4.3152439e-017 lat=0.032395875                lu0=0                          wvth0=1.2499966e-008 wk2=-1.2547231e-009            wcit=-1.3072691e-010            wvoff=-4.0330739e-009 weta0=1.152e-007                 wetab=1.4688e-008                wua=8.9676591e-017 wub=2.6812127e-026             wuc=8.9283068e-018             wa0=3.7628459e-007 wags=3.9656308e-008             wketa=-2.1325396e-009            wpclm=-1.47712e-008 wpdiblc2=-1.094e-010                wagidl=1.4576916e-016             wtvoff=-1.58323e-010 wkt1=2.2807112e-009             wua1=1.1059448e-016             wub1=-7.5563636e-026 wuc1=-4.5788364e-018            pvth0=-6.5758889e-015            pk2=2.1646339e-015 pcit=1.4249233e-016             pvoff=1.1750989e-014             pua=1.050432e-022 pub=-1.1183327e-031            puc=-2.9253085e-024            pa0=-7.9544412e-013 pags=1.3961618e-013             pketa=-5.908664e-015             ppclm=-2.0113203e-013 ppdiblc2=1.374926e-015              pagidl=-1.7595683e-022            ptvoff=6.39265e-016 pkt1=1.6168344e-014             pua1=2.153527e-022              pub1=-3.5712364e-031 puc1=-1.0642284e-023            wat=0.0021297332               pat=-1.9188896e-008 wvsat=0                          wu0=2.88e-009                  pu0=0 pvsat=0                          u0_mc=8.25758e-05                lu0_mc=-7.44008e-10 wu0_mc=-2.97273e-11               pu0_mc=2.67843e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.23 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.40147711 k2=-0.0019638134              cit=0.0025840223               voff=-0.17473404 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-2.3847245e-009            ub=3.0942967e-018             uc=5.3452918e-011 vsat=98000                      a0=3.4094686                  ags=1.3700218 keta=-0.097546714               pclm=1.0530667                  pdiblc2=-0.0035688889 agidl=7.4696333e-010             tvoff=0.000470243                kt1=-0.30130308 ute=-1                         ua1=8.9151324e-010             ub1=-7.8444444e-019 uc1=5.2227834e-011             at=307500.29                  lvth0=-4.2631111e-009 lk2=-5.2979549e-009            lcit=-1.7265843e-009            lvoff=-1.4439018e-008 lua=2.7627682e-016             lub=-4.6994987e-025            luc=-2.1446897e-018 la0=-9.0205992e-007            lags=-6.5170654e-007            lketa=6.5056763e-008 lpclm=2.6043733e-007             lpdiblc2=6.2008889e-010             lagidl=-5.2861028e-016 ltvoff=-2.94555e-010              lkt1=2.9987251e-008             lua1=-1.0656848e-016 lub1=3.1004444e-025             luc1=-3.2076339e-017            lat=-0.17589858 lu0=0                          wvth0=4.8184e-009                wk2=1.9110007e-009 wcit=-6.7651201e-010            wvoff=4.6092676e-009             weta0=1.152e-007 wetab=1.4688e-008                wua=2.9366186e-016             wub=-2.0405344e-025 wuc=7.7318451e-018             wa0=-6.5140871e-007            wags=-1.2746144e-007 wketa=1.3949899e-008             wpclm=-1.960192e-007             wpdiblc2=4.352e-010 wagidl=-1.2475576e-016            wtvoff=3.44872e-010               wkt1=3.1181275e-008 wua1=3.3889395e-016             wub1=-3.6224e-025               wuc1=-2.4046416e-017 pvth0=1.7970176e-015             pk2=-1.286005e-015             pcit=7.3739809e-016 pvoff=2.3308367e-015             pua=-1.1730074e-022            pub=1.398102e-031 puc=-1.6211653e-024            pa0=3.2474157e-013             pags=3.2177453e-013 pketa=-2.3438522e-014            ppclm=-3.571712e-015             ppdiblc2=7.81312e-016 pagidl=1.1891534e-022             ptvoff=9.07828e-017               pkt1=-1.533327e-014 pua1=-3.3493729e-023            pub1=-4.46464e-032              puc1=1.0577377e-023 wat=-0.04172036                pat=2.8607705e-008             wvsat=0 wu0=2.88e-009                  pu0=0                          pvsat=0 lvsat=0                          u0_mc=-0.00131111                lu0_mc=7.75107e-10 wu0_mc=4.208e-10                  pu0_mc=-2.23232e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.24 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.37668621 k2=-0.0088550293              cit=-0.0011503126              voff=-0.18279738 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-2.2657003e-009            ub=2.75e-018                  uc=4.960161e-011 vsat=98000                      a0=4.652                      ags=2.1863257 keta=-0.013461155               pclm=1.4756                     pdiblc2=0.00055315936 agidl=-7.7738591e-010            tvoff=0.00048736                 kt1=-0.21043728 ute=-1                         ua1=1.9438707e-011             ub1=1.104e-018 uc1=6.7797899e-011             at=44869.759                  lvth0=1.1603065e-008 lk2=-8.875767e-010             lcit=6.6339003e-010             lvoff=-9.2784757e-009 lua=2.0010133e-016             lub=-2.496e-025                luc=3.2014694e-019 la0=-1.69728e-006              lags=-1.1741411e-006            lketa=1.1242006e-008 lpclm=-9.984e-009                lpdiblc2=-2.018022e-009             lagidl=4.4697323e-016 ltvoff=-3.0551e-010               lkt1=-2.8166861e-008            lua1=4.5155923e-016 lub1=-8.9856e-025               luc1=-4.2041181e-017            lat=-0.0078150459 lu0=0                          wvth0=1.5213348e-008             wk2=1.9031459e-009 wcit=8.7654962e-010             wvoff=3.0447884e-009             weta0=1.152e-007 wetab=1.4688e-008                wua=1.8530229e-016             wub=-5.2992e-026 wuc=7.2087633e-018             wa0=-4.8096e-007               wags=-6.6299847e-007 wketa=-2.602744e-008             wpclm=-1.56672e-007              wpdiblc2=5.2086263e-010 wagidl=2.7167109e-016             wtvoff=3.04312e-010               wkt1=-6.8573952e-009 wua1=5.6414926e-016             wub1=-8.8128e-025               wuc1=-3.2727715e-017 pvth0=-4.8557492e-015            pk2=-1.2809779e-015            pcit=-2.5656135e-016 pvoff=3.3321034e-015             pua=-4.7950612e-023            pub=4.313088e-032 puc=-1.2863929e-024            pa0=2.156544e-013              pags=6.6451823e-013 pketa=2.1469748e-015             ppclm=-2.875392e-014             ppdiblc2=7.2648792e-016 pagidl=-1.3479785e-022            ptvoff=1.16741e-016               pkt1=9.0114785e-015 pua1=-1.7765713e-022            pub1=2.875392e-031              puc1=1.6133409e-023 wat=0.011463092                pat=-5.4297033e-009            wvsat=0 wu0=2.88e-009                  pu0=0                          pvsat=0 lvsat=0                          u0_mc=-0.00088                   lu0_mc=4.992e-10 wu0_mc=2.9664e-10                 pu0_mc=-1.43769e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18_mac.25 nmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.38352036 k2=-0.010941318               cit=-0.00036625255             voff=-0.19906137 eta0=-0.25                      etab=-0.0658                    u0=0.007122449 ua=-1.9391147e-009            ub=1.6838776e-018             uc=3.5876633e-011 vsat=97708.279                  a0=2.5176122                  ags=-3.5611185 keta=0.020332674                pclm=1.6571429                  pdiblc2=-0.018474406 agidl=3.8673953e-010             tvoff=-0.000591918               kt1=-0.3122542 ute=-1.2367347                 ua1=3.9997129e-010             ub1=-6.0816327e-019 uc1=-7.5746939e-011            at=27976.71                   lvth0=8.9377483e-009 lk2=-7.3924006e-011            lcit=3.5760662e-010             lvoff=-2.9355197e-009 lua=7.273293e-017              lub=1.6618776e-025             luc=5.6728883e-018 lvsat=0.00011377115              la0=-8.6486878e-007            lags=1.0673622e-006 lketa=-1.9375876e-009            lpclm=-8.0785714e-008            lpdiblc2=5.4027286e-009 lagidl=-7.0356858e-018            ltvoff=1.15408e-010               lkt1=1.154174e-008 lua1=3.0315152e-016             lub1=-2.3081633e-025            luc1=1.3941306e-017 lat=-0.0012267567              lute=9.2326531e-008             lu0=3.4622449e-009 wvth0=7.6260855e-009             wk2=-2.913439e-009             wcit=4.3335918e-010 wvoff=9.3066741e-009             weta0=1.152e-007                 wetab=1.4688e-008 wua=3.8667833e-017             wub=2.3657143e-025             wuc=1.0485816e-017 wa0=-1.6611722e-007            wags=2.1682809e-006             wketa=-2.0530174e-008 wpclm=-2.8153469e-007            wpdiblc2=6.4339224e-009             wagidl=-9.2412149e-017 wtvoff=6.36204e-010               wkt1=2.1038576e-008             wua1=3.4061178e-016 wub1=-3.9967347e-025            wuc1=1.3139853e-017             pvth0=-1.8967168e-015 pk2=5.974902e-016              pcit=-8.3717082e-017            pvoff=8.89968e-016 pua=9.2368251e-024             pub=-6.9798857e-032            puc=-2.5644433e-024 pa0=9.2865718e-014             pags=-4.3968073e-013            pketa=3.0412359e-018 ppclm=1.9942531e-014             ppdiblc2=-1.5796054e-015            pagidl=7.1946152e-024 ptvoff=-1.26967e-017              pkt1=-1.8679504e-015            pua1=-9.047751e-023 pub1=9.9712653e-032             puc1=-1.7549427e-024            wat=-0.005102529 pat=1.0308886e-009             wvsat=0.00032076222              pvsat=-1.2509727e-010 wu0=4.5844898e-009             pu0=-6.6475102e-016            u0_mc=0.000636738 vsat_mc=1479.59                    lvsat_mc=-0.000577041               lu0_mc=-9.23262e-11 wvsat_mc=-0.000426122               pvsat_mc=1.66188e-10                wu0_mc=-1.14612e-10 pu0_mc=1.66188e-17 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model pch_18_mac.global pmos ( modelid=10                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=0                          igbmod=0 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_18'              permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=3.65e-009                  toxm=3.65e-009                  dtox=4.74e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=1e-008 xw=0                          dlc=1.24e-008                  dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.43 k3=0.2                        k3b=0.4                        w0=0 dvt0=0.5                        dvt1=0.2                        dvt2=-0.09 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.4                       voffl=-5e-009 dvtp0=8e-007                     dvtp1=3                          lpe0=6e-008 lpeb=1e-007                     xj=8.5e-008                   ngate=1.15e+020 ndep=1e+017                     nsd=1e+020                     phin=0.15 cdsc=0                          cdscb=0                          cdscd=0 ud=0                          nfactor=0.8                        a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=1.2 delta=0.02                       pscbe1=9.264e+008                 pscbe2=1e-020 fprout=100                        pdits=0                          pditsd=0 pditsl=0                          rsh=16.7                       rdsw=200 prwg=0                          prwb=0                          wr=1 alpha0=0                          alpha1=0.055                      beta0=13.7 bgidl=9e+008                     cgidl=5                          egidl=0.5 aigbacc=0.01238                    bigbacc=0.006109                   cigbacc=0.2809 nigbacc=4.05                       aigbinv=0.35                       bigbinv=0.03 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1 aigc=0.009898                   bigc=0.001383                   cigc=1.515e-005 aigsd=0.0086                     bigsd=0.0004353                  cigsd=3.925e-020 nigc=1                          poxedge=1                          pigcd=1.672 ntox=1                          cgso=7.5e-012                   cgdo=7.5e-012 cgbo=0                          cgdl=1.105e-010                 cgsl=1.105e-010 clc=0                          cle=0.6                        cf='9.43e-011+5.68e-11*ccoflag_18' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=5                          noff=2.6                        voffcv=-0.092 kt1l=0                          prt=0                          fnoimod=1 tnoimod=1                          em=7.46e+006                  ef=1.15 noia=0                          noib=0                          noic=0 lintnoi=-1.44e-008                 jss=2.81e-07                   jsd=2.81e-07 jsws=4.79e-14                   jswd=4.79e-14                   jswgs=4.79e-14 jswgd=4.79e-14                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=7.34                       bvd=7.34 xjbvs=1                          xjbvd=1                          jtssws=0 jtsswgs=5e-011                     jtsswgd=5e-011                     njtssw=20 njtsswg=8                          xtsswgs=0.46                       xtsswgd=0.46 tnjtsswg=1                          vtsswgs=7                          vtsswgd=7 pbs=0.830                      pbd=0.830                      cjs=0.001836 cjd=0.001836                   mjs=0.451                      mjd=0.451 pbsws=0.924                      pbswd=0.924                      cjsws=1.454e-010 cjswd=1.454e-010                 mjsws=0.560                      mjswd=0.560 pbswgs=0.949                      pbswgd=0.949                      cjswgs=1.847e-010 cjswgd=1.847e-010                 mjswgs=0.678                      mjswgd=0.678 tpb=0.00129                    tcj=0.00085                    tpbsw=0.00107 tcjsw=0.00066                    tpbswg=0.00140                    tcjswg=0.00100 xtis=3                          xtid=3                          dmcg=6.7e-008 dmci=6.7e-008                   dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=-5.1e-009 rshg=14.4                       gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          xrcrg1=12 xrcrg2=1                          pk2we=0                          lk2we=0 wk2we=0                          k2we=0                          pku0we=0 wku0we=-5e-10                     lku0we=0                          ku0we=0 pkvth0we=0                          wkvth0we=0                          lkvth0we=0 kvth0we=-0.005                     wec=-2800                      web=-150 scref=1e-6                       wpemod=1                          rnoia=0 rnoib=0                          tnoia=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.5 sigma_factor='sigma_factor_18' ccoflag='ccoflag_18' rcoflag='rcoflag_18' rgflag='rgflag_18' mismatchflag='mismatchflag_mos_18' globalflag='globalflag_mos_18' totalflag='totalflag_mos_18' global_factor='global_factor_18' local_factor='local_factor_18' sigma_factor_flicker='sigma_factor_flicker_18' noiseflag='noiseflagp_18' noiseflag_mc='noiseflagp_18_mc' delvto=0 mulu0=1 dlc_fmt=2 par1_io='par1_io' par2_io='par2_io' par3_io='par3_io' par4_io='par4_io' par5_io='par5_io' par6_io='par6_io' par7_io='par7_io' par8_io='par8_io' par9_io='par9_io' par10_io='par10_io' par11_io='par11_io' par12_io='par12_io' par13_io='par13_io' par14_io='par14_io' par15_io='par15_io' par16_io='par16_io' par17_io='par17_io' par18_io='par18_io' par19_io='par19_io' par20_io='par20_io' w7_io='2.0857*0.40825' w8_io='0.67082*0.40825' w9_io='0.54772*-0.10446' w10_io='0.54772*0.14211' w11_io='0.54772*-0.14894' w12_io='0.54772*0.78318' tox_c='toxp_18'                  dxl_c='dxlp_18'                  dxw_c='dxwp_18' ddlc_c='ddlcp_18'                 cgo_c='cgop_18'                  cgl_c='cglp_18' cj_c='cjp_18'                   cjsw_c='cjswp_18'                 cjswg_c='cjswgp_18' cf_c='cfp_18'                   dvth_c='dvthp_18'                 dwvth_c='dwvthp_18' dlvth_c='dlvthp_18'                dpvth_c='dpvthp_18'                du0_c='du0p_18' dwu0_c='dwu0p_18'                 dlu0_c='dlu0p_18'                 dpu0_c='dpu0p_18' dk2_c='dk2p_18'                  dwk2_c='dwk2p_18'                 dlk2_c='dlk2p_18' dpk2_c='dpk2p_18'                 dags_c='dagsp_18'                 dwags_c='dwagsp_18' dpdiblc2_c='dpdiblc2p_18'             dlpdiblc2_c='dlpdiblc2p_18'            dvsat_c='dvsatp_18' dwvsat_c='dwvsatp_18'               duc_c='ducp_18'                  dluc_c='dlucp_18' dwuc_c='dwucp_18'                 dpuc_c='dpucp_18'                 dvoff_c='dvoffp_18' dlvoff_c='dlvoffp_18'               dwvoff_c='dwvoffp_18'               dpvoff_c='dpvoffp_18' dpkt1_c='dpkt1p_18'                dltvoff_c='dltvoffp_18'              dkt2_c='dkt2p_18' duc1_c='duc1p_18'                 dlub1_c='dlub1p_18'                dlketa_c='dlketap_18' ss_flag_c='ss_flagp_18'              ff_flag_c='ff_flagp_18'              sf_flag_c='sf_flagp_18' fs_flag_c='fs_flagp_18'              monte_flag_c='monte_flagp_18'          c1f_c='c1fp_18' c2f_c='c2fp_18'                  c3f_c='c3fp_18' global_mc='global_mc_flag_18' tox_g='toxp_18_ms_global'        dxl_g='dxlp_18_ms_global'        dxw_g='dxwp_18_ms_global' cgo_g='cgop_18_ms_global'        cgl_g='cglp_18_ms_global'        cj_g='cjp_18_ms_global' cjsw_g='cjswp_18_ms_global'       cjswg_g='cjswgp_18_ms_global'      cf_g='cfp_18_ms_global' dvth_g='dvthp_18_ms_global'       dwvth_g='dwvthp_18_ms_global'      dlvth_g='dlvthp_18_ms_global' dpvth_g='dpvthp_18_ms_global'      du0_g='du0p_18_ms_global'        dwu0_g='dwu0p_18_ms_global' dlu0_g='dlu0p_18_ms_global'       dpu0_g='dpu0p_18_ms_global'       dk2_g='dk2p_18_ms_global' dwk2_g='dwk2p_18_ms_global'       dlk2_g='dlk2p_18_ms_global'       dpk2_g='dpk2p_18_ms_global' dags_g='dagsp_18_ms_global'       dwags_g='dwagsp_18_ms_global'      dvsat_g='dvsatp_18_ms_global' dwvsat_g='dwvsatp_18_ms_global'     dluc_g='dlucp_18_ms_global'       dlketa_g='dlketap_18_ms_global' ss_flag_g='ss_flagp_18_ms_global'    ff_flag_g='ff_flagp_18_ms_global' monte_flag_g='monte_flagp_18_ms_global'                                        sf_flag_g='sf_flagp_18_ms_global' fs_flag_g='fs_flagp_18_ms_global' weight1=-2.2915882 weight2=1.8541176 weight3=1.0677647 weight4=-0.58823529 weight5=-0.40837059 tox_1=8.0597748e-012 tox_2=-2.813774e-011 tox_3=-2.6572367e-012 tox_4=9.4219297e-011 tox_5=7.1465402e-013 dxl_1=4.8370644e-010 dxl_2=-1.6886243e-009 dxl_3=-1.5947618e-010 dxl_4=-5.6546372e-009 dxl_5=4.2889837e-011 dxl_max=-1.5e-008 dxw_1=-2.1173527e-009 dxw_2=-9.4864039e-010 dxw_3=2.3732503e-010 dxw_4=-3.7265088e-025 dxw_5=-1.1765292e-008 dxw_max=-1.2e-008 cgo_1=-6.0687e-014 cgo_2=3.5716e-014 cgo_3=9.6404e-015 cgo_4=-1.0732e-029 cgo_5=8.2291e-015 cgl_1=-8.9412e-013 cgl_2=5.2622e-013 cgl_3=1.4203e-013 cgl_4=6.9896e-029 cgl_5=1.2124e-013 cj_1=1.4856e-005 cj_2=-8.7433e-006 cj_3=-2.36e-006 cj_4=-1.0173e-021 cj_5=-2.0145e-006 cjsw_1=1.1765e-012 cjsw_2=-6.9242e-013 cjsw_3=-1.8689e-013 cjsw_4=-3.002e-028 cjsw_5=-1.5954e-013 cjswg_1=1.4945e-012 cjswg_2=-8.7957e-013 cjswg_3=-2.3741e-013 cjswg_4=-1.1184e-028 cjswg_5=-2.0266e-013 cf_1=-7.6304e-013 cf_2=4.4907e-013 cf_3=1.2121e-013 cf_4=1.2335e-028 cf_5=1.0347e-013 dvth_1=-0.0058524 dvth_2=-0.0029508 dvth_3=0.00049632 dvth_4=8.846e-019 dvth_5=0.0012874 dwvth_1=-8.4283e-010 dwvth_2=2.6991e-010 dwvth_3=8.6161e-012 dwvth_4=-1.2127e-025 dwvth_5=1.3345e-010 dlvth_1=5.5107e-012 dlvth_2=1.4314e-011 dlvth_3=1.5798e-013 dlvth_4=-5.104e-027 dlvth_5=-2.1038e-012 dpvth_1=-2.2752e-017 dpvth_2=-5.9246e-017 dpvth_3=1.037e-018 dpvth_4=3.3642e-032 dpvth_5=9.0017e-018 du0_1=4.9392e-005 du0_2=0.000151182 du0_3=5.45112e-006 du0_4=-1.18638e-020 du0_5=-2.10762e-005 dwu0_1=2.448595e-011 dwu0_2=4.523955e-011 dwu0_3=5.068635e-012 dwu0_4=-2.385185e-026 dwu0_5=-7.7231e-012 dlu0_1=-1.2014e-013 dlu0_2=5.4883e-014 dlu0_3=6.2137e-012 dlu0_4=4.8332e-028 dlu0_5=1.1889e-013 dpu0_1=1.4019e-018 dpu0_2=7.2864e-019 dpu0_3=-3.0081e-019 dpu0_4=-3.4041e-034 dpu0_5=-3.1086e-019 dk2_1=0.001956 dk2_2=0.0019536 dk2_3=4.0495e-005 dk2_4=5.3353e-019 dk2_5=-0.00049273 dwk2_1=1.1028e-010 dwk2_2=-6.4946e-011 dwk2_3=-5.1324e-013 dwk2_4=-1.4238e-026 dwk2_5=-1.4672e-011 dlk2_1=6.5058e-012 dlk2_2=-3.8103e-012 dlk2_3=-8.3213e-012 dlk2_4=-7.7694e-028 dlk2_5=-1.0029e-012 dpk2_1=4.5083e-017 dpk2_2=1.0373e-017 dpk2_3=-5.8341e-018 dpk2_4=-1.167e-032 dpk2_5=-9.1161e-018 dags_1=0.0013833 dags_2=0.00067001 dags_3=0.0010512 dags_4=4.564e-019 dags_5=-0.00026225 dwags_1=-2.2845e-010 dwags_2=-1.1932e-009 dwags_3=8.2049e-010 dwags_4=4.7756e-025 dwags_5=1.8205e-010 dvsat_1=-503.13 dvsat_2=-851.2 dvsat_3=376 dvsat_4=-7.7169e-013 dvsat_5=183.45 dwvsat_1=1.3657e-005 dwvsat_2=0.00031499 dwvsat_3=0.00023774 dwvsat_4=1.1389e-019 dwvsat_5=-1.8382e-005 dluc_1=1.8332e-019 dluc_2=-1.0882e-019 dluc_3=3.3527e-019 dluc_4=-4.584e-035 dluc_5=-1.8823e-020 dlketa_1=-6.1108e-011 dlketa_2=3.6274e-011 dlketa_3=-1.1176e-010 dlketa_4=-4.4625e-026 dlketa_5=6.2745e-012 ss_flag_1=0.054487 ss_flag_2=-0.031757 ss_flag_3=-0.13012 ss_flag_4=7.1537e-017 ss_flag_5=-0.0094 ff_flag_1=-0.061108 ff_flag_2=0.036274 ff_flag_3=-0.11176 ff_flag_4=-2.9739e-017 ff_flag_5=0.0062745 monte_flag_1=0.0604875 monte_flag_2=-0.211162 monte_flag_3=-0.0199425 monte_flag_4=-0.707113 monte_flag_5=0.00536337 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.9998 b_4=-0.0002176                 c_4=0.0002609                  d_4=-0.001733 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=-0.0025                    mis_a_2=-0.042                     mis_a_3=-0.006 mis_b_1=0.0022                     mis_b_2=-0.1236                    mis_b_3=0.0477 mis_c_1=0.9692                     mis_c_2=0                          mis_c_3=0 mis_d_1=0.0008                     mis_d_2=0                          mis_d_3=0 mis_e_1=0.0051                     mis_e_2=0.0482                     mis_e_3=-0.0277 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=0                          xl0=1e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=60                         co_rsd=16.7                       bidirectionflag=1 designflag=1 cf0=9.43e-011                  cco=5.68e-11 noimod=6                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718                      tnoiamax=1e1 tnoiac1=4162131.0367               tnoiac2=-17357183.454              rnoiamax=0.001 rnoiac1=-0.022218                  rnoiac2=0.74858 saref0=0.468e-6            sbref0=0.468e-6 samax=10e-6               sbmax=10e-6 samin=0.135e-6            sbmin=0.135e-6 rllodflag=0                   lreflod=1e-6                llodref=1 lod_clamp=-1e90 wlod0=0 ku00=-0e-9               lku00=0e-16               wku00=-0e-15 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=-0.6 kvth00=-0e-10              lkvth00=-0.0e-16            wkvth00=-0e-16 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0.0                 lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=-8e-9              lku000=1e-16             wku000=-2.5e-15     		pku000=0 llodku000=1                   wlodku000=1 kvth000=-0e-10             lkvth000=-0.5e-16	      wkvth000=-3.5e-16     		pkvth000=0 llodvth00=1                   wlodvth00=1                  steta000=0 stk200=0.5                 lodk200=1 lodeta000=1 wlod1=0                   llod1=0.4e-6 ku01=-2.35e-7            lku01=15e-14              wku01=1e-14 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=-1 kvth01=0.5e-8              lkvth01=-15e-22             wkvth01=3e-15 pkvth01=0e-29               llodvth1=2                   wlodvth1=1 steta01=1                  lodeta01=1 stk21=-0.0                lodk21=1 wlod2=0 ku02=0                   lku02=0                   wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0 kvth02=0                   lkvth02=0                   wkvth02=0 pkvth02=0                   llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0       		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0                   lku03=0                   wku03=0 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0 kvth03=0                   lkvth03=0                   wkvth03=0 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=0e-2                lku003=-0e-9               wku003=0e-9        		pku003=0 llodku003=1                   wlodku003=1 kvth003=0.000               lkvth003=0.0e-10             wkvth003=0e-9       		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=4.68e-7             sa_b1=1.35e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.98e-7             spamax=16e-7               spamin=1.98e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc='2.0e-6*0'          ldpckvth0='0.6+0.4'           pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc='6.3e-4*0'          ldpcku0='0.5*2'             pku0dpc=0.0e-14 keta0dpc=-0.04               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc='0'                 wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='-0.000'            wkvth0dpl=0                   wdplkvth0=1 lkvth0dpl='-0.5e-7*0'         ldplkvth0='0.8+0.2'           pkvth0dpl=0 ku0dpl='1*0'               wku0dpl=0                   wdplku0=1 lku0dpl='1.70e-3'           ldplku0='0.5'               pku0dpl=-2e-11 keta0dpl=0.05                wketa0dpl=0                   wdplketa0=1 kvsatdpl=0.04                wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=0.0e-6              wkvth0dpx=0                   wdpxkvth0=1 lkvth0dpx=0e-10               ldpxkvth0=1                   pkvth0dpx=0 ku0dpx=0                   wku0dpx=0                   wdpxku0=1 lku0dpx=0                   ldpxku0=1                   pku0dpx=0 keta0dpx=0                   wketa0dpx=0                   wdpxketa0=1 kvsatdpx=0                   wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0.000              wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-10            ldpskvth0=1.0                 pkvth0dps=0 ku0dps=-0.01               wku0dps=0                   wdpsku0=1 lku0dps=0.0e-14             ldpsku0=1                   pku0dps=0 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=0.00                wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa=0.0e-9              ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa=-0.0                wku0dpa=0e-9                wdpaku0=1 lku0dpa=-0e-8               ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                   wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.31e-7             spbmax='16e-7+1.6e-6+0.135e-6'    spbmin='1.98e-7+0.198e-6+0.135e-6' pse_mode=1 kvth0dp2=0.0                 wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=5e-7                ldp2kvth0=0.6                 pkvth0dp2=0 ku0dp2=0.00                wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=2.5e-4              ldp2ku0=0.5                 pku0dp2=0 keta0dp2=-0.00               wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=-0.2                wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.0                wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0e-8               ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=1.0                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=10e-6               enxmax=10e-6		 enxmin=0.18e-6 kvth0enx='-0.025'            wkvth0enx='1e-9'              wenxkvth0=1.0 lkvth0enx='1e-7*0'            lenxkvth0=1.0                 pkvth0enx=-0e-17 ku0enx='-1.20+0.1'         wku0enx='-1.0e-7'           wenxku0=1.0 lku0enx='1e-11'             lenxku0=1.5                 pku0enx='-1.0e-15*0' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx='-0.5*0'            wka0enx=0                   wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx='-1*0'              wenx=0                   ku0enx0='0' eny0=8e-8 enyref=8e-8		 enymax=2.0e-6              enymin=0.045e-6 kvth0eny='-0.005*0'          wkvth0eny='-1.1e-8'           wenykvth0=1 lkvth0eny='1.0e-8*0'          lenykvth0=1.0                 pkvth0eny=0 ku0eny='1.1'               wku0eny='5.0e-7*1.2'        wenyku0=1 ku0eny0='-0.15'             wku0eny0='-1.0e-6*1'         weny0ku0=1 lku0eny='7.8e-7'            lenyku0='1.0'               pku0eny=-0.0e-16 keta0eny='0'                 wketa0eny=-5e-9               wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny='0'                 weny=1e-6 kvth0eny1='(-2.0e-4*0)'      wkvth0eny1='-1.0e-10*0'       weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1='(-8.0e-18)*0' ku0eny1='(-1e-2)*0.3'      wku0eny1='(-1.0e-10)*0'     weny1ku0=1 lku0eny1='(-1.0e-5)*0'      leny1ku0=1.0                pku0eny1='(-5.5e-17)*0' keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1='(1.0e-8)*0'       weny1ka0=1 lka0eny1='(4.0e-9)*0'       leny1ka0=1.0                pka0eny1='(3.0e-15)*0' kvsateny1=-0.0               weny1=1e-6 rx_mode=0 rxref=20e-6           ringxmax=9.027e-6            ringxmin=0.477e-6 kvth0rx='(0.02)*1'          wkvth0rx=-0.0e-5             wrxkvth0=1.0 lkvth0rx='(1.0e-9)*0'        lrxkvth0=1.0                 pkvth0rx=0.0e-17 ku0rx='(1.00)*0.6'        wku0rx=0.0e-4              wrxku0=1.0 lku0rx='(1.0e-5)*0'        lrxku0=1.0                 pku0rx='-1.0e-14*0' keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx='-0.3'              wrx=0                   ku0rx0=0.5 ry_mode=0 ryref=1.008e-5            ringymax=9.027e-6            ringymin=0.477e-6 kvth0ry='0.01*0'            wkvth0ry='-0.0e-5+2e-5*0'    wrykvth0=1.0 lkvth0ry='(1.0e-8)*0'        lrykvth0='1.0+0'             pkvth0ry=0.0e-16 ku0ry='-0.1'              wku0ry='-4.0e-7'           wryku0=1.0 lku0ry='2.5e-5*1'          lryku0='0.8'               pku0ry='(-5.0e-16)*0' keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry='-3.0*0'            wry=1e-6 kvth0ry0='(-0.01)*0'         ku0ry0='-0.09' sfxref=1.89e-7           sfxmax=3e-6               minwodx=0.53e-6 sfxmin=1.89e-7 lrefodx=5e-8              lodxref=1                 wodx=1e-6 kvth0odxa=-0.50             lkvth0odxa=2.0e-13           lodxakvth0=2.0 wkvth0odxa=-1.0e-12          wodxakvth0=2.0               pkvth0odxa=0.0e-16 ku0odxa=4.00              lku0odxa=2.0e-20           lodxaku0=3.0 wku0odxa=-1.0e-12          wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.3 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=0.5               r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.065             lku0odx1a=1.0e-7            lodx1aku0=1.0 wku0odx1a=-1.0e-12          wodx1aku0=2.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-1.5e-4           lkvth0odx1b=0.0e-7            lodx1bkvth0=0.5 wkvth0odx1b=2.0e-16           wodx1bkvth0=2.0               pkvth0odx1b=0.0e-16 ku0odx1b=0.000             lku0odx1b=0.0e-6            lodx1bku0=0.5 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=8.1e-7 sfymin=2.61e-7           sfymax=1e-6              minwody=9e-7 wody=1e-6 kvth0odya=0                 lkvth0odya=0e-5              lodyakvth0=1.0 wkvth0odya=0e-7              wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=-0.5              lku0odya=3.0e-7            lodyaku0=1.0 wku0odya=2.5e-5            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=-0e-2             wketa0ody=0                 wodyketa0=1 kvsatody=-0.0 lrefody=5.0e-8            lodyref=0.5 kvth0odyb=-0.00             lkvth0odyb=3.0e-9            lodybkvth0=1.0 wkvth0odyb=1.0e-8            wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.00             lku0odyb=0.0e-10           lodybku0=1.0 wku0odyb=-0.0e-7           wodybku0=1.0               pku0odyb=-0e-16 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model pch_18_mac.1 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-006                     wmax=0.00090001                 vth0=-0.401958 k2=0.012                      cit=0.001                      voff=-0.14036 eta0=0.01                       etab=-0.04                      u0=0.016 ua=1.79568e-009               ub=1.008e-018                 uc=3.9301875e-011 vsat=100000                     a0=1.9939049                  ags=0.6081735 keta=-0.04                      pclm=0.9                        pdiblc2=0.0009 agidl=4.7253673e-011             tvoff=0.0032832                  kt1=-0.168988 kt2=-0.041                     ute=-0.8                       ua1=3.1290656e-009 ub1=-3.6373047e-018            uc1=5.6e-011                   at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=0                          wk2=0                          wvoff=0 wu0=0                          wuc=0                          wags=0 pvth0=0                          pk2=0                          pvoff=0 pu0=0                          puc=0                          pkt1=0 wvsat=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18_mac.2 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.40115041 k2=0.013223777                cit=0.00092040041              voff=-0.14001767 eta0=0.01                       etab=-0.04                      u0=0.015587121 ua=1.6651222e-009             ub=1.0503889e-018             uc=3.8167749e-011 vsat=100000                     a0=1.987791                   ags=0.57383228 keta=-0.038623737               pclm=0.81742424                 pdiblc2=0.00076237374 agidl=4.2750588e-011             tvoff=0.00322974                 kt1=-0.16566405 kt2=-0.041206439               ute=-0.8                       ua1=3.1444876e-009 ub1=-3.6425649e-018            uc1=5.820202e-011              at=120000 lvth0=-7.2763941e-009            lk2=-1.1026231e-008            lcit=7.171923e-010 lvoff=-3.0843826e-009            lu0=3.7200379e-009             lua=1.1763256e-015 lub=-3.8192389e-025            luc=1.0218479e-017             la0=5.5085825e-008 lags=3.0941442e-007             lketa=-1.2400126e-008            lpclm=7.4400758e-007 lpdiblc2=1.2400126e-009             lagidl=4.0572791e-017             ltvoff=4.81698e-010 lkt1=-2.9948785e-008            lkt2=1.8600189e-009             lua1=-1.3895213e-016 lub1=4.7393878e-026             luc1=-1.9840202e-017            wvth0=0 wk2=0                          wvoff=0                          wu0=0 wuc=0                          wags=0                          pvth0=0 pk2=0                          pvoff=0                          pu0=0 puc=0                          pkt1=0                          wvsat=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18_mac.3 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.40892111 k2=0.011869991                cit=0.0021165083               voff=-0.13438143 eta0=0.01                       etab=-0.04                      u0=0.019 ua=3.2067129e-009             ub=3.4444444e-019             uc=1.5602944e-011 vsat=100000                     a0=1.9381799                  ags=0.56735612 keta=-0.045733333               pclm=1.5                        pdiblc2=0.0024688889 agidl=4.6131159e-011             tvoff=0.00478623                 kt1=-0.17221249 kt2=-0.036093778               ute=-1.0844444                 ua1=2.2689852e-009 ub1=-4.0072544e-018            uc1=-5.5111111e-012            at=134222.22 lvth0=1.1936711e-009             lk2=-9.5506042e-009            lcit=-5.8656533e-010 lvoff=-9.2278838e-009            lu0=0                          lua=-5.0400825e-016 lub=3.8755556e-025             luc=3.4814116e-017             la0=1.0916197e-007 lags=3.1647344e-007             lketa=-4.6506667e-009            lpdiblc2=-6.2008889e-010 lagidl=3.6887969e-017             ltvoff=-1.21488e-009              lkt1=-2.281099e-008 lkt2=-3.7127822e-009            lua1=8.1534545e-016             lub1=4.4490547e-025 luc1=4.9607111e-017             lute=3.1004444e-007             lat=-0.015502222 wvth0=0                          wk2=0                          wvoff=0 wu0=0                          wuc=0                          wags=0 pvth0=0                          pk2=0                          pvoff=0 pu0=0                          puc=0                          pkt1=0 wvsat=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18_mac.4 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-006                     wmax=0.00090001                 vth0=-0.407056 k2=0.0095998443               cit=0.000732                   voff=-0.14001408 eta0=0.01                       etab=-0.04                      u0=0.019 ua=2.9915328e-009             ub=5.56256e-019               uc=2.437e-011 vsat=99809.68                   a0=2.5734947                  ags=0.55202753 keta=-0.0419357                 pclm=1.8588                     pdiblc2=0.00072 agidl=8.4252575e-011             tvoff=0.0034947                  kt1=-0.17739619 kt2=-0.0432912                 ute=-0.6                       ua1=3.779921e-009 ub1=-3.7095711e-018            uc1=5.952e-011                 at=184505.6 lvth0=0                          lk2=-8.0977104e-009            lcit=2.9952e-010 lvoff=-5.6229888e-009            lu0=0                          lua=-3.6629299e-016 lub=2.5199616e-025             luc=2.92032e-017               la0=-2.974395e-007 lags=3.2628373e-007             lketa=-7.081152e-009             lpclm=-2.29632e-007 lpdiblc2=4.992e-010                 lagidl=1.2490263e-017             ltvoff=-3.88303e-010 lkt1=-1.9493422e-008            lkt2=8.93568e-010               lua1=-1.5165344e-016 lub1=2.5438818e-025             luc1=7.9872e-018                lat=-0.047683584 lvsat=0.0001218048               wvth0=0                          wk2=0 wvoff=0                          wu0=0                          wuc=0 wags=0                          pvth0=0                          pk2=0 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18_mac.5 pmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=9e-006                     wmax=0.00090001                 vth0=-0.41077747 k2=-0.00014433861             cit=0.0012040816               voff=-0.16088473 eta0=0.01                       etab=-0.04                      u0=0.018408163 ua=2.711669e-009              ub=7.4692245e-019             uc=4.1122449e-012 vsat=103343.29                  a0=2.7049935                  ags=1.0268346 keta=-0.063106429               pclm=1.6665306                  pdiblc2=0.0014081633 agidl=1.0241774e-010             tvoff=0.00249808                 kt1=-0.20564755 kt2=-0.047510204               ute=-0.6                       ua1=3.661101e-009 ub1=-3.3741003e-018            uc1=1.2261225e-010             at=100859.82 lvth0=1.4513731e-009             lk2=-4.297479e-009             lcit=1.1540816e-010 lvoff=2.5165627e-009             lu0=2.3081633e-010             lua=-2.5714611e-016 lub=1.7763624e-025             luc=3.7103725e-017             la0=-3.4872406e-007 lags=1.4110899e-007             lketa=1.1754321e-009             lpclm=-1.5464694e-007 lpdiblc2=2.3081633e-010             lagidl=5.4058472e-018             ltvoff=3.79455e-013 lkt1=-8.4753888e-009            lkt2=2.5389796e-009             lua1=-1.0531364e-016 lub1=1.2355454e-025             luc1=-1.6618775e-017            lat=-0.01506173 lvsat=-0.0012563031              wvth0=0                          wk2=0 wvoff=0                          wu0=0                          wuc=0 wags=0                          pvth0=0                          pk2=0 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          pvsat=0 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18_mac.6 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-007                     wmax=9e-006                     vth0=-0.402012 k2=0.012074583                cit=0.001                      voff=-0.14063535 eta0=0.01                       etab=-0.04                      u0=0.016222222 ua=1.9158667e-009             ub=9.7666667e-019             uc=3.996e-011 vsat=100000                     a0=1.988877                   ags=0.60761164 keta=-0.040077569               pclm=0.92222222                 pdiblc2=0.00092103125 agidl=4.7240065e-011             tvoff=0.00329244                 kt1=-0.16798667 kt2=-0.041717188               ute=-0.77777778                ua1=3.2659211e-009 ub1=-3.7617004e-018            uc1=6.3111111e-011             at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=4.86e-010                  wk2=-6.7125e-010               wvoff=2.478123e-009 wu0=-2e-009                    wua=-1.08168e-015              wub=2.82e-025 wuc=-5.923125e-018             wa0=4.525035e-008              wags=5.056748e-009 wketa=6.98125e-010               wpclm=-2e-007                    wpdiblc2=-1.8928125e-010 wagidl=1.224697e-019              wtvoff=-8.32e-011                 wkt1=-9.012e-009 wkt2=6.4546875e-009             wute=-2e-007                    wua1=-1.2316996e-015 wub1=1.1195615e-024             wuc1=-6.4e-017                  pvth0=0 pk2=0                          pvoff=0                          pu0=0 puc=0                          pkt1=0                          wvsat=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.7 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-007                     wmax=9e-006                     vth0=-0.40116998 k2=0.013304416                cit=0.00091723845              voff=-0.14030825 eta0=0.01                       etab=-0.04                      u0=0.015811668 ua=1.7837055e-009             ub=1.0220924e-018             uc=3.9027926e-011 vsat=100000                     a0=1.9867391                  ags=0.57366749 keta=-0.038635523               pclm=0.84311771                 pdiblc2=0.00079547452 agidl=4.2736969e-011             tvoff=0.00323612                 kt1=-0.16448258 kt2=-0.041953518               ute=-0.77471942                ua1=3.2933411e-009 ub1=-3.7718775e-018            uc1=6.5988098e-011             at=120000 lvth0=-7.5866452e-009            lk2=-1.1080796e-008            lcit=7.4568159e-010 lvoff=-2.9471485e-009            lu0=3.6990954e-009             lua=1.1907721e-015 lub=-4.0928573e-025            luc=8.3979855e-018             la0=1.9263133e-008 lags=3.0583684e-007             lketa=-1.2992835e-008            lpclm=7.127317e-007 lpdiblc2=1.1312661e-009             lagidl=4.0572898e-017             ltvoff=5.07454e-010 lkt1=-3.1571824e-008            lkt2=2.1293342e-009             lua1=-2.4705421e-016 lub1=9.1694912e-026             luc1=-2.5921654e-017            lute=-2.7555836e-008 wvth0=1.7609318e-010             wk2=-7.257543e-010             wvoff=2.6152048e-009 wu0=-2.0209192e-009            wua=-1.0672495e-015            wub=2.5466852e-025 wuc=-7.741598e-018             wa0=9.4674171e-009             wags=1.4831395e-009 wketa=1.0607402e-010             wpclm=-2.3124116e-007            wpdiblc2=-2.9790708e-010 wagidl=1.2257653e-019             wtvoff=-5.74734e-011              wkt1=-1.0633237e-008 wkt2=6.7237038e-009             wute=-2.2752525e-007            wua1=-1.3396817e-015 wub1=1.1638133e-024             wuc1=-7.0074702e-017            pvth0=2.7922604e-015 pk2=4.9108375e-016             wcit=2.845767e-011              pcit=-2.5640361e-016 pvoff=-1.2351071e-015            pu0=1.8848192e-016             pua=-1.3001859e-022 pub=2.4625659e-031             puc=1.6384442e-023             pa0=3.2240422e-013 pags=3.2198213e-014             pketa=5.3343793e-015             ppclm=2.8148287e-013 ppdiblc2=9.7871872e-016             pagidl=-9.624978e-028             ptvoff=-2.31797e-016 pkt1=1.4607349e-014             pkt2=-2.4238372e-015            pute=2.4800252e-013 pua1=9.7291869e-022             pub1=-3.9870931e-031            puc1=5.4733068e-023 wvsat=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.8 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-007                     wmax=9e-006                     vth0=-0.4099936 k2=0.011710643                cit=0.0021721589               voff=-0.13477664 eta0=0.01                       etab=-0.04                      u0=0.019339338 ua=3.3965975e-009             ub=2.4354437e-019             uc=1.3353216e-011 vsat=100000                     a0=1.8414663                  ags=0.55955418 keta=-0.046783704               pclm=1.4927333                  pdiblc2=0.0025882201 agidl=4.6117898e-011             tvoff=0.00478525                 kt1=-0.17377529 kt2=-0.036745867               ute=-1.0844444                 ua1=2.3578601e-009 ub1=-4.1670581e-018            uc1=-6.8028746e-012            at=135802.47 lvth0=2.0311012e-009             lk2=-9.3435828e-009            lcit=-6.2218169e-010 lvoff=-8.9766048e-009            lu0=-1.4606538e-010            lua=-5.6728016e-016 lub=4.393316e-025              luc=3.6383419e-017             la0=1.7761048e-007 lags=3.2122034e-007             lketa=-4.1113185e-009            lpclm=4.6506667e-009 lpdiblc2=-8.2282663e-010            lagidl=3.6887685e-017             ltvoff=-1.18109e-009 lkt1=-2.1442774e-008            lkt2=-3.5470053e-009            lua1=7.7262003e-016 lub1=5.2244183e-025             luc1=5.3420506e-017             lute=3.1004444e-007 lat=-0.017224691               wvth0=9.65236e-009               wk2=1.4341326e-009 wvoff=3.5568594e-009             wu0=-3.0540444e-009            wua=-1.7089613e-015 wub=9.0810062e-025             wuc=2.0247555e-017             wa0=8.7042228e-007 wags=7.0217399e-008             wketa=9.4533333e-009             wpclm=6.54e-008 wpdiblc2=-1.0739813e-009            wagidl=1.1935323e-019             wtvoff=8.86423e-012 wkt1=1.4065197e-008             wkt2=5.8688e-009                wua1=-7.998745e-016 wub1=1.4382335e-024             wuc1=1.1625871e-017             pvth0=-7.5368704e-015 pk2=-1.863193e-015             wcit=-5.00855e-010              pcit=3.205472e-016 pvoff=-2.2615107e-015            pu0=1.3145884e-015             pua=5.6944721e-022 pub=-4.659844e-031             puc=-1.4123736e-023            pa0=-6.1603658e-013 pags=-4.2722131e-014            pketa=-4.8541333e-015            ppclm=-4.1856e-014 ppdiblc2=1.8246397e-015             pagidl=2.5508907e-027             ptvoff=-3.04105e-016 pkt1=-1.2313945e-014            pkt2=-1.491992e-015             pua1=3.8452884e-022 pub1=-6.9782725e-031            puc1=-3.4320558e-023            wat=-0.014222222 pat=1.5502222e-008             wvsat=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.9 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-007                     wmax=9e-006                     vth0=-0.40656669 k2=0.0099014634               cit=0.000760288                voff=-0.13928838 eta0=0.01                       etab=-0.04                      u0=0.019457778 ua=3.1571022e-009             ub=5.2890667e-019             uc=2.6751244e-011 vsat=98679.2                    a0=2.5804915                  ags=0.52853343 keta=-0.041804796               pclm=1.8986667                  pdiblc2=0.00024920373 agidl=8.4238763e-011             tvoff=0.00363514                 kt1=-0.17590903 kt2=-0.04377744                ute=-0.6                       ua1=3.8757364e-009 ub1=-3.7881719e-018            uc1=7.1125687e-011             at=178152.89 lvth0=-1.6212064e-010            lk2=-8.1857079e-009            lcit=2.8141568e-010 lvoff=-6.0890901e-009            lu0=-2.2186667e-010            lua=-4.140032e-016 lub=2.5669973e-025             luc=2.7808681e-017             la0=-2.9536567e-007 lags=3.4107362e-007             lketa=-7.2978192e-009            lpclm=-2.5514667e-007 lpdiblc2=6.7414388e-010             lagidl=1.2490331e-017             ltvoff=-4.4502e-010 lkt1=-2.0077177e-008            lkt2=9.532016e-010              lua1=-1.9882078e-016 lub1=2.7995466e-025             luc1=3.5462267e-018             lat=-0.04432896 lvsat=0.000845312                wvth0=-4.4038214e-009            wk2=-2.7145717e-009 wvoff=-6.5313e-009               wu0=-4.12e-009                 wua=-1.4901248e-015 wub=2.46144e-025               wuc=-2.14312e-017              wa0=-6.2971622e-008 wags=2.1144694e-007             wketa=-1.1781328e-009            wpclm=-3.588e-007 wpdiblc2=4.2371664e-009             wagidl=1.2430308e-019             wtvoff=-1.26389e-009 wkt1=-1.3384397e-008            wkt2=4.37616e-009               wua1=-8.6233891e-016 wub1=7.0740701e-025             wuc1=-1.0445119e-016            pvth0=1.4590857e-015 pk2=7.9197782e-016             wcit=-2.54592e-010              pcit=1.6293888e-016 pvoff=4.1949114e-015             pu0=1.9968e-015                pua=4.2939187e-022 pub=-4.233216e-032             puc=1.2550668e-023             pa0=-1.8664479e-014 pags=-1.3310903e-013            pketa=1.950005e-015              ppclm=2.29632e-013 ppdiblc2=-1.5744949e-015            pagidl=-6.170112e-028             ptvoff=5.10455e-016 pkt1=5.2537955e-015             pkt2=-5.367024e-016             pua1=4.2450606e-022 pub1=-2.3009831e-031            puc1=3.996876e-023              wat=0.0571744 pat=-3.0191616e-008            wvsat=0.01017432                 pvsat=-6.5115648e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.10 pmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=9e-007                     wmax=9e-006                     vth0=-0.41097908 k2=-0.00021865302             cit=0.0011620644               voff=-0.16155424 eta0=0.01                       etab=-0.04                      u0=0.018560091 ua=2.8051365e-009             ub=7.3100227e-019             uc=3.5260771e-012 vsat=105162.39                  a0=2.7640517                  ags=1.0169229 keta=-0.062722547               pclm=1.6357143                  pdiblc2=0.001392517 agidl=1.0240237e-010             tvoff=0.00248896                 kt1=-0.20512477 kt2=-0.048176446               ute=-0.6                       ua1=3.6664154e-009 ub1=-3.4087997e-018            uc1=1.2887769e-010             at=103169.81 lvth0=1.5587135e-009             lk2=-4.2388625e-009            lcit=1.2472288e-010 lvoff=2.5945967e-009             lu0=1.2823129e-010             lua=-2.7673658e-016 lub=1.7788245e-025             luc=3.6866497e-017             la0=-3.6695417e-007 lags=1.5060174e-007             lketa=8.6010351e-010             lpclm=-1.5259524e-007 lpdiblc2=2.282517e-010              lagidl=5.4065252e-018             ltvoff=1.98752e-012 lkt1=-8.6830372e-009            lkt2=2.6688138e-009             lua1=-1.1718558e-016 lub1=1.319995e-025              luc1=-1.8977054e-017            lat=-0.01508556 lvsat=-0.0016831304              wvth0=1.8145117e-009             wk2=6.6882968e-010 wvoff=6.0256664e-009             wu0=-1.3673469e-009            wua=-8.4120777e-016 wub=1.4328163e-025             wuc=5.2755102e-018             wa0=-5.3152413e-007 wags=8.9205187e-008             wketa=-3.4549346e-009            wpclm=2.7734694e-007 wpdiblc2=1.4081633e-010             wagidl=1.3836739e-019             wtvoff=8.20817e-011 wkt1=-4.7050142e-009            wkt2=5.9961735e-009             wua1=-4.7829612e-017 wub1=3.1229507e-025             wuc1=-5.6389009e-017            pvth0=-9.6606419e-016 pk2=-5.2754874e-016            wcit=3.781551e-010              pcit=-8.383249e-017 pvoff=-7.0230553e-016            pu0=9.2326531e-016             pua=1.7631423e-022 pub=-2.2158367e-033            puc=2.135051e-024              pa0=1.64071e-013 pags=-8.5434752e-014            pketa=2.8379577e-015             ppclm=-1.8465306e-014 ppdiblc2=2.3081633e-017             pagidl=-6.1020912e-027            ptvoff=-1.44725e-017 pkt1=1.868836e-015              pkt2=-1.1685076e-015            pua1=1.0684743e-022 pub1=-7.6004654e-032            puc1=2.122451e-023              wat=-0.020789923 pat=2.1446984e-010             wvsat=-0.016371861               pvsat=3.841446e-009 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.11 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.39531118 k2=0.011410214                cit=0.0009842875               voff=-0.13218809 eta0=-0.05                      etab=-0.04                      u0=0.011 ua=1.479e-010                 ub=1.5e-018                   uc=2.51775e-011 vsat=100000                     a0=1.9452161                  ags=0.59326045 keta=-0.034517813               pclm=1                          pdiblc2=0.00056239688 agidl=4.7282714e-011             tvoff=0.0032                     kt1=-0.184 kt2=-0.036863281               ute=-1                         ua1=8.6057278e-010 ub1=-1.016815e-018             uc1=5.9570313e-011             at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=-5.5447416e-009            wk2=-7.331769e-011             wvoff=-5.1244056e-009 wu0=2.7e-009                   wua=5.0949e-016                wub=-1.89e-025 wuc=7.381125e-018              wa0=8.4545167e-008             wags=1.7972821e-008 wketa=-4.3056562e-009            wpclm=-2.7e-007                  wpdiblc2=1.3348969e-010 wagidl=8.4085695e-020             wkt1=5.4e-009                   wkt2=2.0861719e-009 wua1=9.3311387e-016             wub1=-1.3508354e-024            wuc1=-6.0813281e-017 pvth0=0                          pk2=0                          wcit=1.414125e-011 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          weta0=5.4e-008 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.12 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.39419986 k2=0.012395738                cit=0.00091731156              voff=-0.13117562 eta0=-0.05                      etab=-0.04                      u0=0.010741263 ua=8.7658449e-011             ub=1.4715829e-018             uc=2.0112203e-011 vsat=100000                     a0=1.8757916                  ags=0.55103114 keta=-0.033841827               pclm=0.90125316                 pdiblc2=0.0002957318 agidl=4.2785948e-011             tvoff=0.00307951                 kt1=-0.18575143 kt2=-0.036909975               ute=-1.0275252                 ua1=7.5319206e-010 ub1=-8.7111413e-019            uc1=5.9802496e-011             at=120000 lvth0=-1.0012954e-008            lk2=-8.879572e-009             lcit=6.0345326e-010 lvoff=-9.1224027e-009            lu0=2.3312237e-009             lua=5.4277637e-016 lub=2.5603781e-025             luc=4.5638326e-017             la0=6.2551541e-007 lags=3.8048613e-007             lketa=-6.090632e-009             lpclm=8.8970906e-007 lpdiblc2=2.4026523e-009             lagidl=4.0515864e-017             ltvoff=1.08557e-009 lkt1=1.5780401e-008             lkt2=4.2071303e-010             lua1=9.6750026e-016 lub1=-1.3127651e-024            luc1=-2.0919764e-018            lute=2.4800252e-007 wvth0=-6.09701e-009              wk2=9.2056092e-011             wvoff=-5.6041638e-009 wu0=2.5424455e-009             wua=4.5919282e-016             wub=-1.4987296e-025 wuc=9.2825528e-018             wa0=1.0932018e-007             wags=2.1855857e-008 wketa=-4.208253e-009             wpclm=-2.8356307e-007            wpdiblc2=1.5186137e-010 wagidl=7.84955e-020               wtvoff=8.34744e-011               wkt1=8.5087296e-009 wkt2=2.1845157e-009             wua1=9.4645242e-016             wub1=-1.4468737e-024 wuc1=-6.4507661e-017            pvth0=4.9759387e-015             pk2=-1.4900178e-015 wcit=2.8391873e-011             pcit=-1.2839811e-016            pvoff=4.3226217e-015 pu0=1.4195665e-015             pua=4.5317756e-022             pub=-3.525346e-031 puc=-1.7131864e-023            pa0=-2.2322282e-013            pags=-3.4986149e-014 pketa=-8.7760344e-016            ppclm=1.2220324e-013             ppdiblc2=-1.655289e-016 pagidl=5.0367658e-026             ptvoff=-7.52104e-016              pkt1=-2.8009653e-014 pkt2=-8.8607815e-016            pua1=-1.2018033e-022            pub1=8.653047e-031 puc1=3.3286358e-023             wvsat=0                          weta0=5.4e-008 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.13 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.39996208 k2=0.014883551                cit=0.0020696064               voff=-0.1302703 eta0=-0.13533333                etab=-0.04                      u0=0.0098648889 ua=-1.9077493e-010            ub=2.2490293e-018             uc=4.1381726e-011 vsat=100000                     a0=3.2712492                  ags=0.69613197 keta=-0.028078298               pclm=1.6001667                  pdiblc2=0.0014439355 agidl=4.6047099e-011             tvoff=0.00713096                 kt1=-0.10423673 kt2=-0.028205644               ute=-1.0844444                 ua1=-9.6298657e-010 ub1=1.1255667e-019             uc1=1.402061e-010              at=120000 lvth0=-3.7321336e-009            lk2=-1.1591288e-008            lcit=-6.5254806e-010 lvoff=-1.0109198e-008            lu0=3.2864711e-009             lua=8.4626875e-016 lub=-5.9137877e-025            luc=2.2454545e-017             la0=-8.9553338e-007 lags=2.2232622e-007             lketa=-1.2372878e-008            lpclm=1.2789333e-007 lpdiblc2=1.1511103e-009             lagidl=3.6961209e-017             ltvoff=-3.33051e-009 lkt1=-7.3070624e-008            lkt2=-9.0670076e-009            lua1=2.838135e-015 lub1=-2.3849663e-024            luc1=-8.9731904e-017            lute=3.1004444e-007 wvth0=6.2399706e-010             wk2=-1.4214846e-009            wvoff=-4.9884369e-010 wu0=5.47296e-009               wua=1.5196739e-015             wub=-8.9683584e-025 wuc=-4.9781039e-018            wa0=-4.1638232e-007            wags=-5.270261e-008 wketa=-7.3815313e-009            wpclm=-3.129e-008                wpdiblc2=-4.412519e-011 wagidl=1.8307159e-019             wtvoff=-2.10228e-009              wkt1=-4.8519503e-008 wkt2=-1.8174e-009               wua1=2.1888875e-015             wub1=-2.4134198e-024 wuc1=-1.206822e-016             pvth0=-2.3499591e-015            pk2=1.597416e-016 wcit=-4.0855771e-010            pcit=3.4787694e-016             pvoff=-1.2421772e-015 pu0=-1.7746944e-015            pua=-7.0274682e-022            pub=4.6165494e-031 puc=-1.5877486e-024            pa0=3.4979289e-013             pags=4.628258e-014 pketa=2.58127e-015               ppclm=-1.527744e-013             ppdiblc2=4.8096458e-017 pagidl=-6.3620283e-026            ptvoff=1.63037e-015               pkt1=3.415112e-014 pkt2=3.47601e-015               pua1=-1.4744346e-021            pub1=1.91884e-030 puc1=9.4516611e-023             wvsat=0                          weta0=1.308e-007 leta0=9.3013333e-008             peta0=-8.3712e-014               pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.14 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.40768402 k2=0.0087845904               cit=9.528e-005                 voff=-0.14384124 eta0=0.01                       etab=-0.04                      u0=0.0072 ua=2.0966686e-010             ub=9.74e-019                  uc=-1.17636e-011 vsat=110920                     a0=1.6722643                  ags=0.68710533 keta=-0.031324387               pclm=3.438                      pdiblc2=0.004400916 agidl=8.4356068e-011             tvoff=0.00159134                 kt1=-0.19632062 kt2=-0.04617588                ute=-0.6                       ua1=2.5343215e-009 ub1=-4.2648589e-018            uc1=-1.5456797e-010            at=260554.48 lvth0=1.2099061e-009             lk2=-7.6879531e-009            lcit=6.110208e-010 lvoff=-1.4237958e-009            lu0=4.992e-009                 lua=5.8998601e-016 lub=2.2464e-025                luc=5.6467554e-017             la0=1.2781691e-007 lags=2.2810327e-007             lketa=-1.0295381e-008            lpclm=-1.04832e-006 lpdiblc2=-7.4135725e-010            lagidl=1.2443469e-017             ltvoff=2.14854e-010 lkt1=-1.4136933e-008            lkt2=2.4339432e-009             lua1=5.9985779e-016 lub1=4.1657968e-025             luc1=9.89235e-017               lat=-0.089954865 lvsat=-0.0069888                 wvth0=-3.3982229e-009            wk2=-1.709386e-009 wvoff=-2.4337246e-009            wu0=6.912e-009                 wua=1.162567e-015 wub=-1.5444e-025               wuc=1.323216e-017              wa0=7.5443284e-007 wags=6.8732222e-008             wketa=-1.0610501e-008            wpclm=-1.7442e-006 wpdiblc2=5.0062534e-010             wagidl=1.8728496e-020             wtvoff=5.75533e-010 wkt1=4.9860351e-009             wkt2=6.534756e-009              wua1=3.4493448e-016 wub1=1.1364253e-024             wuc1=9.8673103e-017             pvth0=2.2426171e-016 pk2=3.439985e-016              wcit=3.439152e-010              pcit=-1.3370573e-016 pvoff=-3.8534746e-018            pu0=-2.69568e-015              pua=-4.7419842e-022 pub=-1.34784e-032              puc=-1.3242317e-023            pa0=-3.9952881e-013 pags=-3.1435713e-014            pketa=4.6478106e-015             ppclm=9.43488e-013 ppdiblc2=-3.0054388e-016            pagidl=4.1559299e-026             ptvoff=-8.34321e-017 pkt1=-9.2424084e-017            pkt2=-1.8693698e-015            pua1=-2.9430465e-022 pub1=-3.5306084e-031            puc1=-4.5870786e-023            wat=-0.016987029 pat=1.0871699e-008             wvsat=-0.0008424                 pvsat=5.39136e-010 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.15 pmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.40753894 k2=0.0016329666               cit=0.0015803265               voff=-0.15398485 eta0=0.01                       etab=-0.04                      u0=0.017040816 ua=1.9633418e-009             ub=1.0368184e-018             uc=2.800949e-011 vsat=82890.709                  a0=2.2221681                  ags=1.0038749 keta=-0.072740356               pclm=0.75                       pdiblc2=0.0015826531 agidl=1.023909e-010              tvoff=0.00253363                 kt1=-0.20073526 kt2=-0.045133546               ute=-0.6                       ua1=3.9610468e-009 ub1=-3.4549351e-018            uc1=8.3762173e-011             at=63439.093 lvth0=1.1533251e-009             lk2=-4.8988198e-009            lcit=3.1852653e-011 lvoff=2.5322094e-009             lu0=1.1540816e-009             lua=-9.3947207e-017 lub=2.0014084e-025             luc=4.0956049e-017             la0=-8.6645564e-008 lags=1.0456314e-007             lketa=5.8568467e-009             lpclm=2.5871527e-022 lpdiblc2=3.5776531e-010             lagidl=5.4098825e-018             ltvoff=-1.52639e-010 lkt1=-1.2415225e-008            lkt2=2.0274329e-009             lua1=4.3434947e-017 lub1=1.0070942e-025             luc1=5.9747448e-018             lat=-0.013079865 lvsat=0.0039426237               wvth0=-1.2816169e-009            wk2=-9.9762799e-010 wvoff=-7.8679248e-010            wu0=0                          wua=-8.3592496e-017 wub=-1.3195286e-025            wuc=-1.6759561e-017            wa0=-4.3828852e-008 wags=1.0094838e-007             wketa=5.5610932e-009             wpclm=1.0744898e-006 wpdiblc2=-3.0306122e-011            wagidl=1.4868492e-019             wtvoff=4.18849e-011 wkt1=-8.6555782e-009            wkt2=3.2575638e-009             wua1=-3.1299786e-016 wub1=3.5381694e-025             wuc1=-1.5785043e-017            pvth0=-6.0121464e-016 pk2=6.6412865e-017             wcit=1.7191837e-012             pcit=-2.4928163e-019 pvoff=-6.46157e-016              pu0=0                          pua=1.1803797e-023 pub=-2.2248386e-032            puc=-1.5455461e-024            pa0=-8.8206748e-014 pags=-4.4000015e-014            pketa=-1.6591112e-015            ppclm=-1.5580102e-013 ppdiblc2=-9.3480612e-017            pagidl=-9.1237078e-027            ptvoff=1.24691e-016 pkt1=5.2278051e-015             pkt2=-5.9126487e-016            pua1=-3.7711039e-023 pub1=-4.7843583e-032            puc1=-1.2321092e-024            wat=0.014967725 pat=-1.5906554e-009            wvsat=0.003672648                pvsat=-1.2217327e-009 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.16 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.41310813 k2=0.013181082                cit=0.001031425                voff=-0.1515812 eta0=0.13                       etab=-0.035386                  u0=0.018 ua=1.8686e-009                ub=1.01e-018                  uc=6.053875e-011 vsat=100000                     a0=2.0978593                  ags=0.66021725 keta=-0.05947375                pclm=0.5                        pdiblc2=0.0004288 agidl=4.7195057e-011             tvoff=0.003                      kt1=-0.178 kt2=-0.02799                   ute=-1                         ua1=4.3441234e-009 ub1=-6.1777116e-018            uc1=-1.7997062e-010            at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=4.0656125e-009             wk2=-1.0295863e-009            wvoff=5.3478716e-009 wu0=-1.08e-009                 wua=-4.19688e-016              wub=7.56e-026 wuc=-1.171395e-017             wa0=2.1178692e-009             wags=-1.8183852e-008 wketa=9.17055e-009               wpdiblc2=2.05632e-010               wagidl=1.3142066e-019 wtvoff=1.08e-010                  wkt1=2.16e-009                  wkt2=-2.7054e-009 wua1=-9.4800347e-016            wub1=1.4360488e-024             wuc1=6.8538825e-017 pvth0=0                          pk2=0                          wcit=-1.1313e-011 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          weta0=-4.32e-008 wetab=-2.49156e-009              pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.17 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.41329725 k2=0.014715916                cit=0.00097129289              voff=-0.15207654 eta0=0.13                       etab=-0.035386                  u0=0.01689899 ua=1.5576555e-009             ub=1.1228535e-018             uc=5.9275782e-011 vsat=100000                     a0=1.9711439                  ags=0.6136996 keta=-0.059313123               pclm=0.40366162                 pdiblc2=0.00014374849 agidl=4.2679471e-011             tvoff=0.0030833                  kt1=-0.17124523 kt2=-0.028286997               ute=-1.0275252                 ua1=4.3396751e-009 ub1=-6.4988718e-018            uc1=-2.0025541e-010            at=120000 lvth0=1.7040278e-009             lk2=-1.3828852e-008            lcit=5.4179028e-010 lvoff=4.4630373e-009             lu0=9.920101e-009              lua=2.8016101e-015 lub=-1.0168103e-024            luc=1.1379344e-017             la0=1.1417053e-006 lags=4.1912405e-007             lketa=-1.4472497e-009            lpclm=8.6800884e-007 lpdiblc2=2.5683141e-009             lagidl=4.0685427e-017             ltvoff=-7.50518e-010 lkt1=-6.086044e-008             lkt2=2.6759473e-009             lua1=4.0078882e-017 lub1=2.8936534e-024             luc1=1.827659e-016              lute=2.4800252e-007 wvth0=4.2155827e-009             wk2=-1.1608397e-009            wvoff=5.6823351e-009 wu0=-7.8272727e-010            wua=-3.3460557e-016            wub=3.8440909e-026 wuc=-1.186578e-017             wa0=5.7829898e-008             wags=-1.1985114e-008 wketa=9.546247e-009              wpclm=-1.4863636e-008            wpdiblc2=2.3393236e-010 wagidl=1.3599296e-019             wtvoff=8.14313e-011               wkt1=6.7538284e-010 wkt2=-2.4718923e-009            wua1=-9.9024844e-016            wub1=1.5921155e-024 wuc1=7.5923608e-017             pvth0=-1.3512317e-015            pk2=1.1825935e-015 wcit=-7.5804941e-013            pcit=-9.5100105e-017            pvoff=-3.0135159e-015 pu0=-2.6784273e-015            pua=-7.6659267e-022            pub=3.3480341e-031 puc=1.3679858e-024             pa0=-5.0196538e-013            pags=-5.5850626e-014 pketa=-3.3850299e-015            ppclm=1.3392136e-013             ppdiblc2=-2.5498628e-016 pagidl=-4.1196354e-026            ptvoff=2.39384e-016               pkt1=1.3376401e-014 pkt2=-2.1039046e-015            pua1=3.8062721e-022             pub1=-1.4061613e-030 puc1=-6.6536894e-023            wvsat=0                          weta0=-4.32e-008 wetab=-2.49156e-009              pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.18 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.40721541 k2=0.015032352                cit=0.001980559                voff=-0.13947229 eta0=0.30066667                 etab=-0.035386                  u0=0.028844444 ua=5.6562395e-009             ub=-6.7755556e-019            uc=5.4562239e-011 vsat=100000                     a0=3.4160679                  ags=0.67369554 keta=-0.060365625               pclm=1.6266667                  pdiblc2=0.00091393778 agidl=4.629239e-011              tvoff=0.00221475                 kt1=-0.24681335 kt2=-0.024791644               ute=-1.6533333                 ua1=4.1195056e-009 ub1=-7.1906742e-018            uc1=-3.2069444e-010            at=120000 lvth0=-4.9251831e-009            lk2=-1.4173767e-008            lcit=-5.5830974e-010 lvoff=-9.2756027e-009            lu0=-3.1004444e-009            lua=-1.6658465e-015 lub=9.4563556e-025             luc=1.6517106e-017             la0=-4.3326184e-007 lags=3.5372847e-007             lketa=-3.0002226e-010            lpclm=-4.6506667e-007 lpdiblc2=1.7288078e-009             lagidl=3.6747345e-017             ltvoff=1.962e-010 lkt1=2.1508808e-008             lkt2=-1.1339876e-009            lua1=2.8006367e-016 lub1=3.647718e-024              luc1=3.1404444e-016             lute=9.3013333e-007 wvth0=4.5407943e-009             wk2=-1.501837e-009             wvoff=4.4702273e-009 wu0=-4.776e-009                wua=-1.6377139e-015            wub=6.8352e-025 wuc=-1.209558e-017             wa0=-4.9458445e-007            wags=-4.0586937e-008 wketa=1.0053625e-008             wpclm=-4.56e-008                 wpdiblc2=2.420736e-010 wagidl=5.0614699e-020             wtvoff=5.52474e-010               wkt1=2.8471872e-008 wkt2=-3.66096e-009              wute=3.072e-007                 wua1=-5.5565824e-016 wub1=1.5303248e-024             wuc1=1.2820409e-016             pvth0=-1.7057124e-015 pk2=1.5542806e-015             wcit=-3.6047213e-010            pcit=2.9698824e-016 pvoff=-1.6923184e-015            pu0=1.67424e-015               pua=6.5379541e-022 pub=-3.683328e-031             puc=1.6184687e-024             pa0=1.0016626e-013 pags=-2.4674639e-014            pketa=-3.938072e-015             ppclm=1.67424e-013 ppdiblc2=-2.6386022e-016            pagidl=5.1865946e-026             ptvoff=-2.74052e-016 pkt1=-1.6921773e-014            pkt2=-8.078208e-016             pute=-3.34848e-013 pua1=-9.3076108e-023            pub1=-1.3388095e-030            puc1=-1.2352262e-022 wvsat=0                          weta0=-1.0464e-007               leta0=-1.8602667e-007 peta0=6.69696e-014               wetab=-2.49156e-009              pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.19 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.41941866 k2=0.0039507069               cit=0.0002453415               voff=-0.15237506 eta0=0.01                       etab=-0.035386                  u0=0.024 ua=3.4130052e-009             ub=5.816e-019                 uc=7.3500742e-012 vsat=128080                     a0=4.6720865                  ags=1.1264257 keta=-0.06114159                pclm=-2.376                     pdiblc2=0.010191376 agidl=8.4051888e-011             tvoff=0.00199838                 kt1=-0.18593657 kt2=-0.02099976                ute=0.424                      ua1=6.2035499e-009 ub1=3.4545069e-019             uc1=3.104e-010                 at=188133.19 lvth0=2.8848948e-009             lk2=-7.0815148e-009            lcit=5.5222944e-010 lvoff=-1.0178299e-009            lu0=0                          lua=-2.3017653e-016 lub=1.39776e-025               luc=4.6732891e-017             la0=-1.2371137e-006 lags=6.3981186e-008             lketa=1.9659494e-010             lpclm=2.09664e-006 lpdiblc2=-4.2087528e-009            lagidl=1.2581267e-017             ltvoff=3.34678e-010 lkt1=-1.7452335e-008            lkt2=-3.5607936e-009            lua1=-1.0537247e-015 lub1=-1.1754019e-024            luc1=-8.9856e-017               lute=-3.9936e-007 lat=-0.043605242               lvsat=-0.0179712                 wvth0=2.9384815e-009 wk2=9.0091105e-010             wvoff=2.1745345e-009             wu0=-2.16e-009 wua=-5.6723569e-016            wub=5.7456e-026                wuc=2.9107759e-018 wa0=-8.6547115e-007            wags=-1.6850076e-007            wketa=5.4907883e-009 wpclm=1.39536e-006               wpdiblc2=-2.6262232e-009            wagidl=1.8298604e-019 wtvoff=3.55731e-010               wkt1=-6.2135649e-010            wkt2=-7.0603488e-009 wute=-5.5296e-007               wua1=-1.6364488e-015            wub1=-1.3531419e-024 wuc1=-1.524096e-016             pvth0=-6.802322e-016             pk2=1.6521823e-017 wcit=2.6288199e-010             pcit=-1.0195839e-016            pvoff=-2.2307507e-016 pu0=0                          pua=-3.1310647e-023            pub=3.234816e-032 puc=-7.9855994e-024            pa0=3.3753375e-013             pags=5.719021e-014 pketa=-1.0178564e-015            ppclm=-7.547904e-013             ppdiblc2=1.5718497e-015 pagidl=-3.2851713e-026            ptvoff=-1.48137e-016              pkt1=1.6978935e-015 pkt2=1.367788e-015              pute=2.156544e-013              pua1=5.9862987e-022 pub1=5.0660922e-031             puc1=5.6070144e-023             wat=0.022120465 pat=-1.4157098e-008            wvsat=-0.0101088                 pvsat=6.469632e-009 wetab=-2.49156e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.20 pmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.40677227 k2=-1.8126226e-005            cit=0.0018159699               voff=-0.16317012 eta0=0.01                       etab=-0.035386                  u0=0.017489796 ua=2.6017396e-009             ub=4.5126122e-019             uc=-1.2431551e-011 vsat=76245.946                  a0=2.7601536                  ags=1.0777029 keta=-0.054489395               pclm=4.6038776                  pdiblc2=-0.0035596574 agidl=1.0247858e-010             tvoff=0.00227369                 kt1=-0.2406208 kt2=-0.030018735               ute=-0.6                       ua1=3.7405818e-009 ub1=-2.5025679e-018            uc1=8.9469388e-011             at=99311.004 lvth0=-2.0471942e-009            lk2=-5.5336699e-009            lcit=-6.0315635e-011 lvoff=3.1922466e-009             lu0=2.5389796e-009             lua=8.6217053e-017 lub=1.9060812e-025             luc=5.4447725e-017             la0=-4.9145989e-007 lags=8.2983086e-008             lketa=-2.3977611e-009            lpclm=-6.2551225e-007 lpdiblc2=1.1541503e-009             lagidl=5.3948564e-018             ltvoff=2.27305e-010 lkt1=3.8745159e-009             lkt2=-4.3393469e-011            lua1=-9.3167113e-017 lub1=-6.4674649e-026            luc1=-3.6930612e-018            lat=-0.0089645894 lvsat=0.002244081                wvth0=-1.695616e-009             wk2=-1.0603785e-010 wvoff=4.1732576e-009             wu0=-2.4244898e-010            wua=-4.2832734e-016 wub=1.84248e-025               wuc=5.0786008e-018             wa0=-3.34341e-007 wags=6.1081273e-008             wketa=-4.2944258e-009            wpclm=-1.0066041e-006 wpdiblc2=2.7465415e-009             wagidl=1.0133957e-019             wtvoff=1.82248e-010 wkt1=1.2882614e-008             wkt2=-4.9044343e-009            wua1=-1.9394678e-016 wub1=-1.6046134e-025            wuc1=-1.8866939e-017            pvth0=1.1270658e-015 pk2=4.092319e-016              wcit=-1.2552823e-010            pcit=4.9521594e-017 pvoff=-1.0025771e-015            pu0=-7.478449e-016             pua=-8.5484904e-023 pub=-1.710072e-032             puc=-8.8310511e-024            pa0=1.3039299e-013 pags=-3.2346785e-014            pketa=2.798377e-015              ppclm=1.8197559e-013 ppdiblc2=-5.2352852e-016            pagidl=-1.0095906e-027            ptvoff=-8.04784e-017 pkt1=-3.568655e-015             pkt2=5.2698137e-016             pua1=3.6054074e-023 pub1=4.1463814e-032             puc1=3.9885061e-024             wat=-0.0044031077 pat=-3.8129044e-009            wvsat=0.0072608197               pvsat=-3.045197e-010 wetab=-2.49156e-009 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.21 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.4072178 k2=0.010337252                cit=0.001                      voff=-0.1493905 eta0=0.01                       etab=-0.031111                  u0=0.011 ua=-1.868576e-010             ub=1.58e-018                  uc=1.5755e-011 vsat=100000                     a0=2.3196728                  ags=0.61152644 keta=-0.041525                  pclm=-1.1                       pdiblc2=0.00124 agidl=4.7193824e-011             tvoff=0.0026812                  kt1=-0.196 kt2=-0.041175                  ute=-1                         ua1=7.1821e-010 ub1=-1.0431195e-018            uc1=3.944625e-011              at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=1.9450944e-009             wk2=-5.80752e-012              wvoff=4.55922e-009 wu0=1.44e-009                  wua=3.2027674e-016             wub=-1.296e-025 wuc=4.4082e-018                wa0=-7.7735002e-008            wags=-6.5515968e-010 wketa=2.709e-009                 wpclm=5.76e-007                  wpdiblc2=-8.64e-011 wagidl=1.3186454e-019             wtvoff=2.22769e-010               wkt1=8.64e-009 wkt2=2.0412e-009                wua1=3.5732536e-016             wub1=-4.1240438e-025 wuc1=-1.045125e-017             pvth0=0                          pk2=0 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          wetab=-4.03056e-009 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.22 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.40853166 k2=0.011188961                cit=0.00097321277              voff=-0.15093456 eta0=0.01                       etab=-0.031111                  u0=0.010724748 ua=-3.0922078e-010            ub=1.6391793e-018             uc=1.6069992e-011 vsat=100000                     a0=2.2673298                  ags=0.56836068 keta=-0.042595044               pclm=-1.4578283                 pdiblc2=0.00094503939 agidl=4.2691464e-011             tvoff=0.00260815                 kt1=-0.19710407 kt2=-0.042413292               ute=-1.0275252                 ua1=5.4311156e-010 ub1=-7.9594151e-019            uc1=4.8032709e-011             at=120000 lvth0=1.1837875e-008             lk2=-7.6738936e-009            lcit=2.4135296e-010 lvoff=1.3911999e-008             lu0=2.4800252e-009             lua=1.1024922e-015 lub=-5.3320543e-025            luc=-2.8380789e-018            la0=4.7161053e-007 lags=3.8892346e-007             lketa=9.6410982e-009             lpclm=3.2240328e-006 lpdiblc2=2.6575951e-009             lagidl=4.0566257e-017             ltvoff=6.58202e-010 lkt1=9.9476913e-009             lkt2=1.1157014e-008             lua1=1.5776369e-015 lub1=-2.2270741e-024            luc1=-7.7364e-017               lute=2.4800252e-007 wvth0=2.4999686e-009             wk2=1.0886413e-010             wvoff=5.2712225e-009 wu0=1.44e-009                  wua=3.3746988e-016             wub=-1.4743636e-025 wuc=3.6883045e-018             wa0=-4.8797016e-008            wags=4.3368952e-009 wketa=3.5277386e-009             wpclm=6.5527273e-007             wpdiblc2=-5.4532364e-011 wagidl=1.3167534e-019             wtvoff=2.52486e-010               wkt1=9.9845646e-009 wkt2=2.6135739e-009             wua1=3.7651445e-016             wub1=-4.6093941e-025 wuc1=-1.3460115e-017            pvth0=-4.9994166e-015            pk2=-1.0331916e-015 wcit=-1.4492045e-012            pcit=1.3057333e-017             pvoff=-6.4151422e-015 pu0=-2.7655242e-029            pua=-1.5491023e-022            pub=1.6070564e-031 puc=6.486258e-024              pa0=-2.6073125e-013            pags=-4.4978415e-014 pketa=-7.3768351e-015            ppclm=-7.1424727e-013            ppdiblc2=-2.871274e-016 pagidl=1.7047297e-027             ptvoff=-2.67755e-016              pkt1=-1.2114527e-014 pkt2=-5.1570885e-015            pua1=-1.7289368e-022            pub1=4.3730063e-031 puc1=2.7109869e-023             wvsat=0                          wetab=-4.03056e-009 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.23 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.38154078 k2=0.011988572                cit=0.00093172194              voff=-0.12962813 eta0=0.01                       etab=-0.031111                  u0=0.0058888889 ua=-6.134567e-010             ub=1.3512729e-018             uc=-5.636298e-011 vsat=100000                     a0=3.98                       ags=1.1020547 keta=-0.030066444               pclm=1.5                        pdiblc2=0.0034844622 agidl=4.6059707e-011             tvoff=0.00312333                 kt1=-0.18733668 kt2=-0.038709056               ute=-0.8                       ua1=1.493459e-009 ub1=-3.1315556e-018            uc1=1.2949345e-010             at=120000 lvth0=-1.758218e-008             lk2=-8.5454701e-009            lcit=2.8657796e-010 lvoff=-9.3120175e-009            lu0=7.7511111e-009             lua=1.4341094e-015 lub=-2.1938745e-025            luc=7.6113861e-017             la0=-1.3952e-006 lags=-1.92803e-007              lketa=-4.0150756e-009            lpdiblc2=-1.1037582e-010 lagidl=3.6894873e-017             ltvoff=9.66513e-011               lkt1=-6.9876267e-010 lkt2=7.1193956e-009             lua1=5.4175819e-016             lub1=3.1874522e-025 luc1=-1.6615621e-016            wvth0=-4.702071e-009             wk2=-4.0607631e-010 wvoff=9.2632973e-010             wu0=3.488e-009                 wua=6.1937674e-016 wub=-4.685824e-026             wuc=2.7837498e-017             wa0=-6.976e-007 wags=-1.9479623e-007            wketa=-8.5408e-010               wpdiblc2=-6.833152e-010 wagidl=1.3438066e-019             wtvoff=2.25386e-010               wkt1=7.060272e-009 wkt2=1.349308e-009              wua1=3.8971854e-016             wub1=6.904214e-026 wuc1=-3.3863555e-017            pvth0=2.8508066e-015             pk2=-4.7190649e-016 wcit=1.71092e-011               pcit=-7.171328e-018             pvoff=-1.6792091e-015 pu0=-2.23232e-015              pua=-4.6218871e-022            pub=5.1075482e-032 puc=-1.9836363e-023            pa0=4.46464e-013               pags=1.7207669e-013 pketa=-2.6006528e-015            ppdiblc2=3.9824589e-016             pagidl=-1.2440719e-027 ptvoff=-2.38215e-016              pkt1=-8.9270477e-015            pkt2=-3.7790387e-015 pua1=-1.8728613e-022            pub1=-1.4037926e-031            puc1=4.9349619e-023 wvsat=0                          wetab=-4.03056e-009              pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.24 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.41019377 k2=0.0030112652               cit=0.0010100272               voff=-0.13574839 eta0=0.01                       etab=-0.031111                  u0=0.02424 ua=3.8688396e-009             ub=-1.794912e-019             uc=-4.4396586e-011 vsat=100000                     a0=2.6424                     ags=0.16970637 keta=-0.01205236                pclm=1.5                        pdiblc2=0.0039535594 agidl=8.4189551e-011             tvoff=0.00425066                 kt1=-0.20644631 kt2=-0.034075087               ute=-2.36                      ua1=-2.307265e-009 ub1=-3.8165232e-018            uc1=-5.702416e-010             at=247972.97 lvth0=7.557289e-010              lk2=-2.7999937e-009            lcit=2.3646256e-010 lvoff=-5.3950491e-009            lu0=-3.9936e-009               lua=-1.4345603e-015 lub=7.6030157e-025             luc=6.8455368e-017             la0=-5.39136e-007 lags=4.0389992e-007             lketa=-1.554409e-008             lpdiblc2=-4.1059799e-010 lagidl=1.2491773e-017             ltvoff=-6.24839e-010              lkt1=1.1531397e-008 lkt2=4.1536559e-009             lua1=2.9742215e-015             lub1=7.5712446e-025 luc1=2.8167422e-016             lute=9.984e-007                 lat=-0.081902698 wvth0=-3.8247875e-010            wk2=1.2391101e-009             wvoff=-3.8110656e-009 wu0=-2.2464e-009               wua=-7.3133609e-016            wub=3.3144883e-025 wuc=2.1539574e-017             wa0=-1.34784e-007              wags=1.7591819e-007 wketa=-1.2181334e-008            wpdiblc2=-3.806091e-010             wagidl=1.3342746e-019 wtvoff=-4.55089e-010              wkt1=6.7621511e-009             wkt2=-2.353231e-009 wute=4.4928e-007                wua1=1.4274445e-015             wub1=1.4516871e-025 wuc1=1.6462138e-016             pvth0=8.6267511e-017             pk2=-1.5248258e-015 wcit=-1.2404879e-011            pcit=1.1717683e-017             pvoff=1.3527238e-015 pu0=1.437696e-015              pua=4.022675e-022              pub=-1.9104104e-031 puc=-1.5805691e-023            pa0=8.626176e-014              pags=-6.5180536e-014 pketa=4.64879e-015               ppdiblc2=2.0451398e-016             pagidl=-6.3402394e-028 ptvoff=1.97289e-016               pkt1=-8.7362503e-015            pkt2=-1.4094138e-015 pute=-2.875392e-013             pua1=-8.5143076e-022            pub1=-1.8910027e-031 puc1=-7.7680737e-023            wat=0.00057814631              pat=-3.7001364e-010 wvsat=0                          wetab=-4.03056e-009              pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18_mac.25 pmos ( level=54                         lmin=1.35e-07                   lmax=3.8e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.43056114 k2=0.0092244197               cit=0.0014678742               voff=-0.17816288 eta0=0.01                       etab=-0.031111                  u0=0.015183674 ua=1.0447253e-009             ub=9.8960408e-019             uc=9.0370204e-011 vsat=64593.959                  a0=-0.66702041                ags=1.4452466 keta=-0.082719775               pclm=1.855102                   pdiblc2=0.00059302106 agidl=1.0240033e-010             tvoff=0.000713536                kt1=-0.18769954 kt2=-0.015727666               ute=0.67346939                 ua1=6.4417772e-009 ub1=-1.6708538e-018            uc1=1.4050524e-010             at=192818.71 lvth0=8.6990057e-009             lk2=-5.223124e-009             lcit=5.7902235e-011 lvoff=1.1146601e-008             lu0=-4.6163265e-010            lua=-3.3315567e-016 lub=3.0435441e-025             luc=1.589632e-017              la0=7.5153796e-007 lags=-9.3560752e-008            lketa=1.2016202e-008             lpclm=-1.384898e-007 lpdiblc2=9.0001195e-010             lagidl=5.3895702e-018             ltvoff=7.54639e-010 lkt1=4.2201587e-009             lkt2=-3.0018384e-009            lua1=-4.3790491e-016 lub1=-7.9686595e-026            luc1=4.4829561e-018             lute=-1.8465306e-007 lat=-0.06039254                lvsat=0.013808356                wvth0=6.8683768e-009 wk2=-3.4333544e-009            wvoff=9.5706487e-009             wu0=5.877551e-010 wua=1.3219782e-016             wub=-9.5554286e-027            wuc=-3.1930031e-017 wa0=8.9944163e-007             wags=-7.1234461e-008            wketa=5.8685113e-009 wpclm=-1.7044898e-008            wpdiblc2=1.2515773e-009             wagidl=1.2951093e-019 wtvoff=7.43905e-010               wkt1=-6.1690383e-009            wkt2=-1.0049219e-008 wute=-4.5844898e-007            wua1=-1.1663771e-015            wub1=-4.5987843e-025 wuc1=-3.7239846e-017            pvth0=-2.7415662e-015            pk2=2.9743537e-016 wcit=-2.1379709e-013            pcit=6.9631606e-018             pvoff=-3.8661447e-015 pu0=3.3237551e-016             pua=6.5489276e-023             pub=-5.8049383e-032 puc=5.0474545e-024             pa0=-3.1708624e-013            pags=3.1208997e-014 pketa=-2.3906498e-015            ppclm=6.6475102e-015             ppdiblc2=-4.3203871e-016 pagidl=8.9342537e-028             ptvoff=-2.70319e-016              pkt1=-3.6930865e-015 pkt2=1.5920216e-015             pute=6.6475102e-014             pua1=1.6015968e-022 pub1=4.6868114e-032             puc1=1.0451399e-024             wat=-0.038065883 pat=1.4701158e-008             wvsat=0.011455535                pvsat=-4.4676587e-009 wetab=-4.03056e-009 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_18ud15_mac.global nmos ( modelid=11                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=0                          igbmod=0 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_18ud15'          permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=3.36e-009                  toxm=3.36e-009                  dtox=2.83e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=1e-008 xw=0                          dlc=1.17e-008                  dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.31 k3=-5.1                       k3b=0.25                       w0=0 dvt0=0.0103                     dvt1=0.02                       dvt2=-0.09 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.4                       voffl=-5e-009 dvtp0=1.5e-006                   dvtp1=0                          lpe0=8e-008 lpeb=5e-009                     xj=6.7e-008                   ngate=4.8e+020 ndep=1e+017                     nsd=1e+020                     phin=0.15 cdsc=0                          cdscb=0                          cdscd=0 ud=0                          nfactor=0.7                        a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=0.45 delta=0.01                       pscbe1=9.264e+008                 pscbe2=1e-020 fprout=750                        pdits=0                          pditsd=0 pditsl=0                          rsh=18.0                       rdsw=150 prwg=0                          prwb=0                          wr=1 alpha0=0                          alpha1=0.06                       beta0=8.83 bgidl=1.1e+009                   cgidl=5                          egidl=0.8 aigbacc=0.01238                    bigbacc=0.006109                   cigbacc=0.2809 nigbacc=4.05                       aigbinv=0.35                       bigbinv=0.03 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1 aigc=0.009898                   bigc=0.001383                   cigc=1.515e-005 aigsd=0.0086                     bigsd=0.0004353                  cigsd=3.925e-020 nigc=1                          poxedge=1                          pigcd=1.672 ntox=1                          cgso=4.5e-011                   cgdo=4.5e-011 cgbo=0                          cgdl=7.9e-011                   cgsl=7.9e-011 clc=0                          cle=0.6                        cf='8.09e-011+5.742e-11*ccoflag_18ud15' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=5                          noff=3                          voffcv=-0.085 kt1l=0                          prt=0                          fnoimod=1 tnoimod=1                          em=2.53e+009                  ef=0.94 noia=0                          noib=0                          noic=0 lintnoi=-3.80e-008                 jss=2.69e-07                   jsd=2.69e-07 jsws=7.06e-14                   jswd=7.06e-14                   jswgs=7.06e-14 jswgd=7.06e-14                   njs=1.09                       njd=1.09 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=7.9                        bvd=7.9 xjbvs=1                          xjbvd=1                          jtsswgs=2e-009 jtsswgd=2e-009                     njtsswg=15                         xtsswgs=0.5 xtsswgd=0.5                        tnjtsswg=1                          vtsswgs=1 vtsswgd=1                          pbs=0.715                      pbd=0.715 cjs=0.001472                   cjd=0.001472                   mjs=0.336 mjd=0.336                      pbsws=0.457                      pbswd=0.457 cjsws=1.086e-010                 cjswd=1.086e-010                 mjsws=0.015 mjswd=0.015                      pbswgs=0.923                      pbswgd=0.923 cjswgs=2.016e-010                 cjswgd=2.016e-010                 mjswgs=0.552 mjswgd=0.552                      tpb=0.00137                    tcj=0.00079 tpbsw=0.00230                    tcjsw=0.00020                    tpbswg=0.00114 tcjswg=0.00073                    xtis=3                          xtid=3 dmcg=6.7e-008                   dmci=6.7e-008                   dmdg=0 dmcgt=0                          dwj=0                          xgw=0 xgl=2.64e-009                  rshg=16.42                      gbmin=1e-012 rbpb=50                         rbpd=50                         rbps=50 rbdb=50                         rbsb=50                         ngcon=1 xrcrg1=12                         xrcrg2=1                          pk2we=0 lk2we=0                          wk2we=0                          k2we=0 pku0we=-1e-16                     wku0we=0                          lku0we=0 ku0we=-0.004                     pkvth0we=-1e-17                     wkvth0we=0 lkvth0we=0                          kvth0we=0.0085                     wec=-2800 web=-150                       scref=1e-6                       wpemod=1 rnoia=0                          rnoib=0                          tnoia=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.5 sigma_factor='sigma_factor_18ud15' ccoflag='ccoflag_18ud15' rcoflag='rcoflag_18ud15' rgflag='rgflag_18ud15' mismatchflag='mismatchflag_mos_18ud15' globalflag='globalflag_mos_18ud15' totalflag='totalflag_mos_18ud15' global_factor='global_factor_18ud15' local_factor='local_factor_18ud15' sigma_factor_flicker='sigma_factor_flicker_18ud15' noiseflag='noiseflagn_18ud15' noiseflag_mc='noiseflagn_18ud15_mc' delvto=0 mulu0=1 dlc_fmt=2 par1_io='par1_io' par2_io='par2_io' par3_io='par3_io' par4_io='par4_io' par5_io='par5_io' par6_io='par6_io' par7_io='par7_io' par8_io='par8_io' par9_io='par9_io' par10_io='par10_io' par11_io='par11_io' par12_io='par12_io' par13_io='par13_io' par14_io='par14_io' par15_io='par15_io' par16_io='par16_io' par17_io='par17_io' par18_io='par18_io' par19_io='par19_io' par20_io='par20_io' w1_io='2.0857*0.40825' w2_io='0.67082*-0.40825' w3_io='0.54772*0.26807' w4_io='0.54772*-0.6902' w5_io='0.54772*-0.32981' w6_io='0.54772*0.098267' tox_c='toxn_18ud15'              dxl_c='dxln_18ud15'              dxw_c='dxwn_18ud15' ddlc_c='ddlcn_18ud15'             cgo_c='cgon_18ud15'              cgl_c='cgln_18ud15' cj_c='cjn_18ud15'               cjsw_c='cjswn_18ud15'             cjswg_c='cjswgn_18ud15' cf_c='cfn_18ud15'               dvth_c='dvthn_18ud15'             dwvth_c='dwvthn_18ud15' dlvth_c='dlvthn_18ud15'            dpvth_c='dpvthn_18ud15'            du0_c='du0n_18ud15' dwu0_c='dwu0n_18ud15'             dlu0_c='dlu0n_18ud15'             dpu0_c='dpu0n_18ud15' dk2_c='dk2n_18ud15'              dwk2_c='dwk2n_18ud15'             dlk2_c='dlk2n_18ud15' dpk2_c='dpk2n_18ud15'             dags_c='dagsn_18ud15'             dwags_c='dwagsn_18ud15' dpdiblc2_c='dpdiblc2n_18ud15'         dlpdiblc2_c='dlpdiblc2n_18ud15'        dvsat_c='dvsatn_18ud15' dwvsat_c='dwvsatn_18ud15'           duc_c='ducn_18ud15'              dluc_c='dlucn_18ud15' dwuc_c='dwucn_18ud15'             dpuc_c='dpucn_18ud15'             dketa_c='dketan_18ud15' dlketa_c='dlketan_18ud15'           dwketa_c='dwketan_18ud15'           dpketa_c='dpketan_18ud15' monte_flag_c='monte_flagn_18ud15'      c1f_c='c1fn_18ud15'              c2f_c='c2fn_18ud15' c3f_c='c3fn_18ud15' global_mc='global_mc_flag_18ud15' tox_g='toxn_18ud15_ms_global'    dxl_g='dxln_18ud15_ms_global' dxw_g='dxwn_18ud15_ms_global'    cgo_g='cgon_18ud15_ms_global' cgl_g='cgln_18ud15_ms_global'    cj_g='cjn_18ud15_ms_global' cjsw_g='cjswn_18ud15_ms_global'   cjswg_g='cjswgn_18ud15_ms_global' cf_g='cfn_18ud15_ms_global'     dvth_g='dvthn_18ud15_ms_global' dwvth_g='dwvthn_18ud15_ms_global'  dlvth_g='dlvthn_18ud15_ms_global' dpvth_g='dpvthn_18ud15_ms_global'  du0_g='du0n_18ud15_ms_global' dwu0_g='dwu0n_18ud15_ms_global'   dlu0_g='dlu0n_18ud15_ms_global' dpu0_g='dpu0n_18ud15_ms_global'   dk2_g='dk2n_18ud15_ms_global' dwk2_g='dwk2n_18ud15_ms_global'   dlk2_g='dlk2n_18ud15_ms_global' dpk2_g='dpk2n_18ud15_ms_global'   dags_g='dagsn_18ud15_ms_global' dwags_g='dwagsn_18ud15_ms_global'  dvsat_g='dvsatn_18ud15_ms_global' dwvsat_g='dwvsatn_18ud15_ms_global' dluc_g='dlucn_18ud15_ms_global' dlketa_g='dlketan_18ud15_ms_global' monte_flag_g='monte_flagn_18ud15_ms_global' weight1=2.2047059 weight2=-1.8575882 weight3=-0.90158824 weight4=-0.58823529 weight5=-0.40471765 tox_1=-2.3955414e-011 tox_2=-8.9373236e-012 tox_3=-1.6291481e-012 tox_4=9.4219297e-011 tox_5=5.1583358e-013 dxl_1=-1.4376247e-009 dxl_2=-5.3637536e-010 dxl_3=-9.7773875e-011 dxl_4=-5.6546372e-009 dxl_5=3.0957612e-011 dxl_max=-2.2e-008 dxw_1=7.0729697e-010 dxw_2=-2.6725306e-009 dxw_3=-7.8365641e-010 dxw_4=4.2997794e-025 dxw_5=-1.1643341e-008 dxw_max=-1.2e-008 cgo_1=3.7272e-013 cgo_2=-2.2768e-013 cgo_3=-6.1739e-014 cgo_4=-2.8927e-029 cgo_5=7.9899e-014 cgl_1=6.5432e-013 cgl_2=-3.9971e-013 cgl_3=-1.0839e-013 cgl_4=-2.848e-029 cgl_5=1.4027e-013 cj_1=-1.2192e-005 cj_2=7.4477e-006 cj_3=2.0195e-006 cj_4=7.2531e-022 cj_5=-2.6136e-006 cjsw_1=-8.9949e-013 cjsw_2=5.4947e-013 cjsw_3=1.49e-013 cjsw_4=3.1935e-029 cjsw_5=-1.9282e-013 cjswg_1=-1.6698e-012 cjswg_2=1.02e-012 cjswg_3=2.7659e-013 cjswg_4=5.9716e-029 cjswg_5=-3.5795e-013 cf_1=6.7006e-013 cf_2=-4.0932e-013 cf_3=-1.1099e-013 cf_4=-1.9574e-029 cf_5=1.4364e-013 dvth_1=-0.0017428 dvth_2=0.008148 dvth_3=0.0018262 dvth_4=-3.0783e-019 dvth_5=-0.0020616 dwvth_1=-6.5967e-010 dwvth_2=7.2666e-010 dwvth_3=6.096e-011 dwvth_4=-9.2199e-027 dwvth_5=-2.0574e-010 dlvth_1=-2.158761e-010 dlvth_2=3.345166e-010 dlvth_3=8.974691e-011 dlvth_4=3.283335e-028 dlvth_5=-9.395166e-011 dpvth_1=4.6949e-017 dpvth_2=4.1044e-017 dpvth_3=2.2304e-017 dpvth_4=-1.1223e-032 dpvth_5=-6.5162e-018 du0_1=0.00015496 du0_2=0.00028363 du0_3=5.1554e-005 du0_4=-2.3503e-021 du0_5=-5.9431e-005 dwu0_1=7.763e-011 dwu0_2=9.4157e-011 dwu0_3=-6.7442e-012 dwu0_4=-6.9556e-027 dwu0_5=-1.6664e-011 dlu0_1=2.1018e-011 dlu0_2=2.2904e-011 dlu0_3=-1.9334e-012 dlu0_4=-2.8615e-027 dlu0_5=-3.5708e-012 dpu0_1=1.1718e-017 dpu0_2=5.39912e-018 dpu0_3=-8.6297e-019 dpu0_4=3.7638e-034 dpu0_5=-9.3827e-019 dk2_1=0.0004774 dk2_2=0.00094815 dk2_3=0.00018641 dk2_4=-7.4278e-020 dk2_5=-0.00019284 dwk2_1=-7.3502e-012 dwk2_2=3.9212e-012 dwk2_3=1.1925e-011 dwk2_4=4.8506e-028 dwk2_5=-2.2095e-012 dlk2_1=3.3952e-011 dlk2_2=7.7131e-011 dlk2_3=1.2768e-011 dlk2_4=-1.1238e-026 dlk2_5=-1.6938e-011 dpk2_1=-4.101e-018 dpk2_2=2.8935e-018 dpk2_3=-6.6306e-018 dpk2_4=-8.8094e-034 dpk2_5=-4.4646e-019 dags_1=0.0021372 dags_2=0.0029623 dags_3=-0.0027687 dags_4=5.229e-019 dags_5=-0.00038734 dwags_1=-2.9389e-009 dwags_2=-1.1743e-009 dwags_3=-6.8702e-010 dwags_4=6.9762e-025 dwags_5=7.139e-011 dvsat_1=51.986 dvsat_2=-15.831 dvsat_3=-308.43 dvsat_4=-1.1821e-014 dvsat_5=28.89 dwvsat_1=7.4621e-005 dwvsat_2=3.73695e-005 dwvsat_3=-4.2311e-005 dwvsat_4=1.1036e-020 dwvsat_5=-1.6368e-005 dluc_1=-1.7928e-019 dluc_2=1.3227e-019 dluc_3=-3.9862e-019 dluc_4=3.9001e-035 dluc_5=-1.3081e-020 dlketa_1=8.9641e-011 dlketa_2=-6.6135e-011 dlketa_3=1.9931e-010 dlketa_4=-1.4829e-026 dlketa_5=6.5405e-012 monte_flag_1=-0.179775 monte_flag_2=-0.0670738 monte_flag_3=-0.0122266 monte_flag_4=-0.707113 monte_flag_5=0.00387125 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.9998 b_4=-0.0009597                 c_4=-0.00141                   d_4=-0.001335 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.0035                     mis_a_2=-0.0405                    mis_a_3=0.0339 mis_b_1=0.001                      mis_b_2=0                          mis_b_3=0 mis_c_1=0.5                        mis_c_2=0                          mis_c_3=0 mis_d_1=0.00087                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.0061                     mis_e_2=-0.076                     mis_e_3=0.0329 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=0                          xl0=1e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0                       bidirectionflag=1 designflag=1 cf0=8.09e-011                  cco=5.742e-11 noimod=6                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718                      tnoiamax=9593223.1145 tnoiac1=123552.3055                tnoiac2=9231959.0635               rnoiamax=0.61424 rnoiac1=0.0085845                  rnoiac2=0.58914 saref0=0.468e-6            sbref0=0.468e-6 samax=10e-6               sbmax=10e-6 samin=0.135e-6            sbmin=0.135e-6 rllodflag=0                   lreflod=1e-6                llodref=1 lod_clamp=-1e90 wlod0=0 ku00=0e-9                lku00=0e-15               wku00=0e-15 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=0 kvth00=-0e-10            lkvth00=-0e-16              wkvth00=-0e-16 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                 lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=3e-9                lku000=1e-15               wku000=1e-15       		pku000=0 llodku000=1                   wlodku000=1 kvth000=-2.5e-10              lkvth000=-3e-16            wkvth000=-6e-16     		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0.2                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=-1e-7               lku01=-1.5e-14            wku01=2e-14 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0.2 kvth01=2e-8                lkvth01=3e-22               wkvth01=3e-15 pkvth01=4.5e-29             llodvth1=2                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=-0.15               lodk21=1 wlod2=0 ku02=0                   lku02=0                   wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0 kvth02=0                   lkvth02=0                   wkvth02=0 pkvth02=0                   llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0                   lku03=0                   wku03=0 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0 kvth03=0                   lkvth03=0                   wkvth03=0 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=0                   lku003=0                   wku003=0         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=4.68e-7             sa_b1=1.35e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.98e-7             spamax=1.6e-6              spamin=1.98e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=0.01                wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl=0.8e-10             ldplkvth0=1.36                pkvth0dpl=0.0e-19 ku0dpl=0.0                 wku0dpl=0e-8                wdplku0=1 lku0dpl=3.2e-6              ldplku0=0.8                 pku0dpl=0.0e-11 keta0dpl=0.5                 wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0.5                 wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx=-0.0                wku0dpx=0e-9                wdpxku0=1 lku0dpx=0.0e-8              ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=0.00                wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps=0.0                 wku0dps=-0.0e-9             wdpsku0=1 lku0dps=0.0e-16             ldpsku0=1.0                 pku0dps=0.0e-23 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=-0.00               wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa=0.0e-9              ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa=0.00                wku0dpa=0e-7                wdpaku0=1 lku0dpa=0.0e-11             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=-0.0                wka0dpa=0                   wdpaka0=1 lka0dpa=-0.0e-7             ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=1.0                 wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.31e-7             spbmax='1.6e-6+1.6e-6+0.135e-6'    spbmin='1.98e-7+1.98e-7+0.135e-6' pse_mode=1 kvth0dp2=0.004               wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0.7e-8              ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.000               wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=0.35e-5             ldp2ku0=0.7                 pku0dp2=0 keta0dp2=0.1                 wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0.8                 wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=1.0                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=10e-6               enxmax=10e-6		 enxmin=0.18e-6 kvth0enx='0.010*3'           wkvth0enx='0.7e-8*2'          wenxkvth0=1 lkvth0enx='4e-5*0'            lenxkvth0=1.0                 pkvth0enx=-3.3e-16 ku0enx='-0.60-0.2'         wku0enx='-0.8e-7*1'         wenxku0=1 lku0enx='0.2e-7'            lenxku0=1                   pku0enx=-3.7e-15 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx='0.0-1'             wka0enx=0                   wenxka0=1 lka0enx='1.0e-7*0'          lenxka0=1.0                 pka0enx='1.0e-14*0' kvsatenx='0.65*1'            wenx=0                   ku0enx0='0.10' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.045e-6 kvth0eny='0.01'              wkvth0eny='3.5e-8*1'          wenykvth0=1 lkvth0eny='1e-7*0'            lenykvth0=1.0                 pkvth0eny=0 ku0eny='(-0.5)*1'          wku0eny='(-0.2e-7)*1'       wenyku0=1 ku0eny0='0.41+0.01'         wku0eny0='-1e-7*2'           weny0ku0=1 lku0eny='(1.2e-11)*1'       lenyku0='1.5'               pku0eny='5.0e-19*0' keta0eny=0.00                wketa0eny=0                   wenyketa0=1 ka0eny='-0.50*1'           wka0eny='-2e-7*0'           wenyka0=1 lka0eny='-6.0e-8*0'         lenyka0=1.0                 pka0eny='(1.0e-14)*0' kvsateny='-0.6+0.4'          weny=1e-6 kvth0eny1=0.000              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=0 ku0eny1='(0.15)*0'         wku0eny1=0.0e-8             weny1ku0=1 lku0eny1='0.0e-5'           leny1ku0=1.0                pku0eny1=-0.0e-14 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1.0                pka0eny1=0 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=2e-5	         ringxmax=9.027e-6		 ringxmin=4.770e-07 kvth0rx=-0.1                wkvth0rx=-1.0e-8             wrxkvth0=1.0 lkvth0rx=0.0e-9              lrxkvth0=1.0                 pkvth0rx=0.0e-16 ku0rx=1.00                wku0rx=1.0e-8              wrxku0=1.0 lku0rx='1.0e-7'            lrxku0=1.0                 pku0rx=0.0e-15 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.0                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=12e-6               ringymax=9.027e-6		 ringymin=0.477e-6 kvth0ry='-0.005'            wkvth0ry='-1e-8*5'           wrykvth0=1.0 lkvth0ry=0.0e-8              lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry=0.1                 wku0ry='1.0e-7*0.3'        wryku0=1.0 lku0ry='1e-5*1'            lryku0=1                   pku0ry=-0.0e-16 keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry=0.0                 wry=1e-6 kvth0ry0=-0.00               ku0ry0=0.01 sfxref=1.89e-7           sfxmax=3e-6               minwodx=0.53e-6 sfxmin=0.189e-6 lrefodx=5e-8              lodxref=1                 wodx=1e-6 kvth0odxa=-0.200            lkvth0odxa=1.0e-13           lodxakvth0=2.0 wkvth0odxa=1.0e-11           wodxakvth0=2.0               pkvth0odxa=0.0e-16 ku0odxa=-0.30             lku0odxa=3.0e-13           lodxaku0=2.0 wku0odxa=5.0e-11           wodxaku0=2.0               pku0odxa=-0.0e-26 keta0odx=0.10              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0005           lkvth0odx1b=0.0e-7            lodx1bkvth0=0.5 wkvth0odx1b=-0.0e-15          wodx1bkvth0=2.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.001            lku0odx1b=0.0e-7            lodx1bku0=0.5 wku0odx1b=-0.5e-14          wodx1bku0=2.0               pku0odx1b=0.0e-16 sfyref=8.1e-7 sfymin=0.15e-6 sfymax=3e-6              minwody=0e-7              wody=1e-6 kvth0odya=-0.000            lkvth0odya=1.0e-13           lodyakvth0=2.0 wkvth0odya=0.0e-6            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=-2.00             lku0odya=2.0e-13           lodyaku0=2.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=0.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.00             lkvth0odyb=-3.0e-9           lodybkvth0=1.0 wkvth0odyb=-7.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=0.10              lku0odyb=0.0e-9            lodybku0=0.8 wku0odyb=-0.0e-5           wodybku0=1.0               pku0odyb=0.0e-13 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_18ud15_mac.1 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-006                     wmax=0.00090001                 vth0=0.43516 k2=0.014574632                cit=0.0015                     voff=-0.17146719 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.5470274e-009            ub=2.510615e-018              uc=1.01528e-010 vsat=100000                     a0=1.8                        ags=0.77816907 keta=-0.060714323               pclm=0.2365                     pdiblc2=0.001 agidl=4.7909339e-010             tvoff=0.001815                   kt1=-0.198016 kt2=-0.03                      ute=-1                         ua1=2.2203714e-009 ub1=-2.08e-018                 uc1=-3.5e-011                  at=120000 lvth0=0                          lk2=0                          luc=0 lketa=0                          lpdiblc2=0                          lu0=0 wvth0=0                          wk2=0                          wuc=0 wags=0                          wketa=0                          pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18ud15_mac.2 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-006                     wmax=0.00090001                 vth0=0.43583426 k2=0.01610097                 cit=0.0015550505               voff=-0.17176577 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.5479495e-009            ub=2.5120759e-018             uc=1.0290646e-010 vsat=100275.25                  a0=1.8421412                  ags=0.71539931 keta=-0.058904163               pclm=0.17959154                 pdiblc2=0.0009583364 agidl=5.1730707e-010             tvoff=0.00183644                 kt1=-0.19457754 kt2=-0.03                      ute=-1                         ua1=2.2881347e-009 ub1=-2.1212879e-018            uc1=-3.6238636e-011            at=121126.33 lvth0=-6.0750761e-009            lk2=-1.3752307e-008            lcit=-4.9600505e-010 lvoff=2.6902347e-009             lua=8.3079606e-018             lub=-1.3162734e-026 luc=-1.2419966e-017            lvsat=-0.0024800252              la0=-3.7969187e-007 lags=5.6555552e-007             lketa=-1.6309534e-008            lpclm=5.1274522e-007 lpdiblc2=3.7538902e-010             lagidl=-3.4430524e-016            ltvoff=-1.93194e-010 lkt1=-3.0980476e-008            lua1=-6.1054678e-016            lub1=3.7200379e-025 luc1=1.1160114e-017             lat=-0.010148263               lu0=0 wvth0=0                          wk2=0                          wuc=0 wags=0                          wketa=0                          pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18ud15_mac.3 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-006                     wmax=0.00090001                 vth0=0.42963686 k2=0.0074962214               cit=0.0011                     voff=-0.16750235 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.4981584e-009            ub=2.5566613e-018             uc=9.36624e-011 vsat=98000                      a0=1.7875156                  ags=0.80265184 keta=-0.064214382               pclm=0.65                       pdiblc2=0.00031105711 agidl=2.9517105e-010             tvoff=0.0017434                  kt1=-0.2102 kt2=-0.03                      ute=-1                         ua1=1.641984e-009 ub1=-1.5524444e-018            uc1=-1.32e-011                 at=194043.2 lvth0=6.8009024e-010             lk2=-4.3731311e-009            lvoff=-1.9568951e-009 lua=-4.5964306e-017            lub=-6.1760853e-026            luc=-2.343936e-018 la0=-3.2014996e-007            lags=4.7045026e-007             lketa=-1.0521396e-008 lpdiblc2=1.0809234e-009             lagidl=-1.0217698e-016            ltvoff=-9.17732e-011 lkt1=-1.3952e-008               lua1=9.375744e-017              lub1=-2.4803556e-025 luc1=-1.3952e-017               lat=-0.089627648               lu0=0 wvth0=0                          wk2=0                          wuc=0 wags=0                          wketa=0                          pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18ud15_mac.4 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-006                     wmax=0.00090001                 vth0=0.43995888 k2=0.0052985221               cit=0.000944                   voff=-0.1757704 eta0=0.18                       etab=-0.035                     u0=0.024 ua=-1.6427414e-009            ub=2.6595534e-018             uc=9.2652e-011 vsat=98503.496                  a0=2.6980475                  ags=0.66058977 keta=-0.1215324                 pclm=0.728                      pdiblc2=-0.00018914922 agidl=1.2975302e-010             tvoff=0.00173603                 kt1=-0.21162952 kt2=-0.03                      ute=-0.688                     ua1=2.7247733e-009 ub1=-2.4704e-018               uc1=-3.5e-011                  at=97009.2 lvth0=-5.9260032e-009            lk2=-2.9666036e-009            lcit=9.984e-011 lvoff=3.334656e-009              lua=4.656883e-017              lub=-1.2761174e-025 luc=-1.69728e-018              lvsat=-0.00032223759             la0=-9.0289038e-007 lags=5.6136999e-007             lketa=2.6162136e-008             lpclm=-4.992e-008 lpdiblc2=1.4010555e-009             lagidl=3.6905546e-018             ltvoff=-8.70605e-011 lkt1=-1.3037107e-008            lua1=-5.992277e-016             lub1=3.39456e-025 lat=-0.027525888               lute=-1.9968e-007               lu0=0 wvth0=0                          wk2=0                          wuc=0 wags=0                          wketa=0                          pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18ud15_mac.5 nmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=9e-006                     wmax=0.00090001                 vth0=0.42400175 k2=-0.0041934273              cit=0.00084489796              voff=-0.17859039 eta0=0.18                       etab=-0.035                     u0=0.019857143 ua=-1.6888162e-009            ub=2.2035268e-018             uc=8.137551e-011 vsat=99853.575                  a0=1.5873206                  ags=2.277551 keta=-0.056962347               pclm=0.68877551                 pdiblc2=0.0042338257 agidl=6.1972392e-011             tvoff=0.00101524                 kt1=-0.25633722 kt2=-0.03                      ute=-1.2                       ua1=1.5469318e-009 ub1=-1.777551e-018             uc1=-4.9795918e-011            at=25175.832 lvth0=2.9727943e-010             lk2=7.3525667e-010             lcit=1.384898e-010 lvoff=4.4344523e-009             lua=6.4537988e-017             lub=5.0238616e-026 luc=2.700551e-018              lvsat=-0.00084876841             la0=-4.6970691e-007 lags=-6.9244898e-008            lketa=9.7981531e-010             lpclm=-3.4622449e-008 lpdiblc2=-3.2390473e-010            lagidl=3.0125e-017                ltvoff=1.94047e-010 lkt1=4.3988975e-009             lua1=-1.3986951e-016            lub1=6.9244898e-026 luc1=5.7704082e-018             lat=0.00048912553              lu0=1.6157143e-009 wvth0=0                          wk2=0                          wuc=0 wags=0                          wketa=0                          pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18ud15_mac.6 nmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=9e-006                     wmax=0.00090001                 vth0=0.38283784 k2=0.0015154251               cit=-6.1728395e-006            voff=-0.16864467 pvoff=0                          wvoff=0                          eta0=0.18 etab=-0.035                     u0=0.031                      ua=-1.1176729e-009 ub=1.7759259e-018             uc=2.0222938e-010             vsat=95894.108 a0=6.4153927                  ags=3.8641975                  keta=-0.15394383 pclm=1.0434568                  pdiblc2=0.0032901235               agidl=9.3990116e-010 tvoff=0.00255089                 kt1=-0.24204914                kt2=-0.055802469 ute=-2.7481482                 ua1=-2.4002254e-010            ub1=-3.5706173e-018 uc1=-2.2158025e-010            at=17737.85                   lvth0=6.2660459e-009 lk2=-9.2526926e-011            lcit=2.6189506e-010             lvoff=2.9923236e-009 lua=-1.8277795e-017            lub=1.1224074e-025             luc=-1.482326e-017 lvsat=-0.00027464561             la0=-1.1697773e-006            lags=-2.9930864e-007 lketa=1.504213e-008              lpclm=-8.6051235e-008            lpdiblc2=-1.870679e-010 lagidl=-9.7174671e-017            ltvoff=-2.86214e-011              lkt1=2.3271247e-009 lua1=1.1923887e-016             lub1=3.2923951e-025             luc1=3.0679136e-017 lat=0.001567633                lute=2.2448148e-007             lu0=0 lkt2=3.741358e-009              wvth0=0                          wk2=0 wuc=0                          wags=0                          wketa=0 pvth0=0                          pk2=0                          puc=0 pketa=0                          wvsat=0                          wu0=0 pu0=0                          pvsat=0                          voff_mc=-0.00516049 pvoff_mc=0.0                        wvoff_mc=0.0                        lvoff_mc=7.48272e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_18ud15_mac.7 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-007                     wmax=9e-006                     vth0=0.43536861 k2=0.014923896                cit=0.0015362917               voff=-0.17107143 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.5469007e-009            ub=2.5162389e-018             uc=1.0250889e-010 vsat=100000                     a0=1.7667745                  ags=0.77929598 keta=-0.061386044               pclm=0.23777778                 pdiblc2=0.00099777778 agidl=4.8625058e-010             tvoff=0.00184031                 kt1=-0.19767822 kt2=-0.03                      ute=-1                         ua1=2.229546e-009 ub1=-2.0944444e-018            uc1=-3.625e-011                at=120000 lvth0=0                          lk2=0                          luc=0 lketa=0                          lpdiblc2=0                          lu0=0 wvth0=-1.8775e-009               wk2=-3.1433799e-009            wcit=-3.26625e-010 wvoff=-3.56181e-009              weta0=-1.6e-007                  wetab=-5e-009 wua=-1.1406e-018               wub=-5.0615e-026               wuc=-8.828e-018 wa0=2.9902927e-007             wags=-1.0142204e-008            wketa=6.04549e-009 wpclm=-1.15e-008                 wpdiblc2=2e-011                     wagidl=-6.4414719e-017 wtvoff=-2.278e-010                wkt1=-3.04e-009                 wua1=-8.257142e-017 wub1=1.3e-025                   wuc1=1.125e-017                 pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.8 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-007                     wmax=9e-006                     vth0=0.43590596 k2=0.01649581                 cit=0.001597866                voff=-0.17133744 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.5483953e-009            ub=2.5176355e-018             uc=1.0396895e-010 vsat=100275.25                  a0=1.8060001                  ags=0.71664671 keta=-0.059691733               pclm=0.1787514                  pdiblc2=0.00095758632 agidl=5.253547e-010              tvoff=0.00186195                 kt1=-0.19437984 kt2=-0.03                      ute=-1                         ua1=2.2996729e-009 ub1=-2.1387907e-018            uc1=-3.7721836e-011            at=121089.39 lvth0=-4.8414984e-009            lk2=-1.4162942e-008            lcit=-5.5478509e-010 lvoff=2.3967598e-009             lua=1.3466952e-017             lub=-1.2583373e-026 luc=-1.3155156e-017            lvsat=-0.0024800252              la0=-3.5342229e-007 lags=5.6446997e-007             lketa=-1.526574e-008             lpclm=5.3182764e-007 lpdiblc2=3.6212502e-010             lagidl=-3.5232809e-016            ltvoff=-1.94944e-010 lkt1=-2.9718418e-008            lua1=-6.318435e-016             lub1=3.9955962e-025 luc1=1.3261246e-017             lat=-0.0098153888              lu0=0 wvth0=-6.4529147e-010            wk2=-3.5535595e-009            wcit=-3.853398e-010 wvoff=-3.8549592e-009            weta0=-1.6e-007                  wetab=-5e-009 wua=4.0126654e-018             wub=-5.0036282e-026            wuc=-9.5623737e-018 wa0=3.2526969e-007             wags=-1.1226547e-008            wketa=7.0881252e-009 wpclm=7.5612374e-009             wpdiblc2=6.7507197e-012             wagidl=-7.242866e-017 wtvoff=-2.29548e-010              wkt1=-1.7793434e-009            wua1=-1.0384451e-016 wub1=1.5752525e-025             wuc1=1.3348801e-017             pvth0=-1.1102199e-014 pk2=3.6957182e-015             pcit=5.2902039e-016             pvoff=2.641274e-015 pua=-4.6430921e-023            pub=-5.2142531e-033            puc=6.6167074e-024 pa0=-2.3642619e-013            pags=9.769928e-015              pketa=-9.3941432e-015 ppclm=-1.7174175e-013            ppdiblc2=1.1937602e-016             pagidl=7.220561e-023 ptvoff=1.57482e-017               pkt1=-1.1358516e-014            pua1=1.9167051e-022 pub1=-2.4800252e-031            puc1=-1.8910193e-023            wat=0.00033250505 pat=-2.9958705e-009            wvsat=0                          wu0=0 pu0=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.9 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-007                     wmax=9e-006                     vth0=0.43133578 k2=0.0069306501               cit=0.0010730864               voff=-0.16930915 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.485957e-009             ub=2.5603284e-018             uc=9.2971407e-011 vsat=98000                      a0=1.7524593                  ags=0.78149618 keta=-0.061446508               pclm=0.71407407                 pdiblc2=0.00013786191 agidl=2.9400029e-010             tvoff=0.0017208                  kt1=-0.20691654 kt2=-0.03                      ute=-1                         ua1=1.6023032e-009 ub1=-1.495679e-018             uc1=-1.0385185e-011            at=192442.77 lvth0=1.3999437e-010             lk2=-3.7369182e-009            lcit=1.7224691e-011 lvoff=1.8592332e-010             lua=-5.4590802e-017            lub=-5.9118586e-026 luc=-1.1678341e-018            la0=-2.9506285e-007            lags=4.9378405e-007 lketa=-1.3353035e-008            lpclm=-5.1674074e-008            lpdiblc2=1.2556246e-009 lagidl=-1.0015178e-016            ltvoff=-4.10981e-011              lkt1=-1.6053412e-008 lua1=1.282895e-016              lub1=-3.014321e-025             luc1=-1.6535704e-017 lat=-0.08759057                lu0=0                          wvth0=-1.5290302e-008 wk2=5.090142e-009              wcit=2.4222222e-010             wvoff=1.6261224e-008 weta0=-1.6e-007                  wetab=-5e-009                    wua=-1.0981246e-016 wub=-3.3003111e-026            wuc=6.2189333e-018             wa0=3.1550616e-007 wags=1.9040097e-007             wketa=-2.4910859e-008            wpclm=-5.7666667e-007 wpdiblc2=1.5587568e-009             wagidl=1.0536865e-017             wtvoff=2.03318e-010 wkt1=-2.9551111e-008            wua1=3.5712711e-016             wub1=-5.1088889e-025 wuc1=-2.5333333e-017            pvth0=4.8608628e-015             pk2=-5.7259164e-015 pcit=-1.5502222e-016            pvoff=-1.9285366e-014            pua=7.7638462e-023 pub=-2.3780409e-032            puc=-1.0584917e-023            pa0=-2.2578395e-013 pags=-2.1000406e-013            pketa=2.548475e-014              ppclm=4.6506667e-013 ppdiblc2=-1.5723107e-015            pagidl=-1.8226812e-023            ptvoff=-4.56075e-016 pkt1=1.8912711e-014             pua1=-3.1078855e-022            pub1=4.8056889e-031 puc1=2.3253333e-023             wat=0.014403911                pat=-1.8333703e-008 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.10 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-007                     wmax=9e-006                     vth0=0.4417723 k2=0.0054507845               cit=0.00096133333              voff=-0.17468974 eta0=0.19777778                 etab=-0.034444444               u0=0.024 ua=-1.6498193e-009            ub=2.6739037e-018             uc=9.3575283e-011 vsat=98559.44                   a0=2.787875                   ags=0.63581794 keta=-0.12567426                pclm=0.70266667                 pdiblc2=-3.6296727e-006 agidl=1.3617223e-010             tvoff=0.00183725                 kt1=-0.20953947 kt2=-0.03                      ute=-0.65333333                ua1=2.7936121e-009 ub1=-2.5144e-018               uc1=-3.3795556e-011            at=99058.349 lvth0=-6.5393762e-009            lk2=-2.7898043e-009            lcit=8.8746667e-011 lvoff=3.629499e-009              lua=5.0281044e-017             lub=-1.3180683e-025 luc=-1.5543147e-018            lvsat=-0.00035804177             la0=-9.5772887e-007 lags=5.8701812e-007             lketa=2.7752725e-008             lpclm=-4.4373333e-008 lpdiblc2=1.3461792e-009             lagidl=8.5817738e-019             ltvoff=-1.15626e-010 lkt1=-1.4374741e-008            lua1=-6.3414818e-016            lub1=3.5054933e-025 luc1=-1.5530667e-018            lat=-0.027824544               lute=-2.2186667e-007 lu0=0                          wvth0=-1.6320762e-008            wk2=-1.3703621e-009 wcit=-1.56e-010                 wvoff=-9.7259296e-009            weta0=-1.6e-007 wetab=-5e-009                    wua=6.3700638e-017             wub=-1.2915335e-025 wuc=-8.30955e-018              wa0=-8.0844748e-007            wags=2.2294652e-007 wketa=3.7276713e-008             wpclm=2.28e-007                  wpdiblc2=-1.6696759e-009 wagidl=-5.7772834e-017            wtvoff=-9.11e-010                 wkt1=-1.881048e-008 wua1=-6.1954928e-016            wub1=3.96e-025                  wuc1=-1.084e-017 pvth0=5.5203573e-015             pk2=-1.5911938e-015            pcit=9.984e-017 pvoff=-2.6535875e-015            pua=-3.3409919e-023            pub=3.7755744e-032 puc=-1.286688e-024             pa0=4.9354638e-013             pags=-2.3083321e-013 pketa=-1.4315296e-014            ppclm=-4.992e-014                ppdiblc2=4.938863e-016 pagidl=2.5491395e-023             ptvoff=2.57088e-016               pkt1=1.2038707e-014 pua1=3.1428434e-022             pub1=-9.984e-032                puc1=1.39776e-023 wat=-0.018442343               pat=2.6878995e-009             wvsat=-0.00050349624 pvsat=3.2223759e-010             wute=-3.12e-007                 pute=1.9968e-013 wu0=0                          pu0=0                          u0_mc=3.46667e-05 lu0_mc=-2.21867e-11               wu0_mc=-3.12e-10                  pu0_mc=1.9968e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.11 nmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=9e-007                     wmax=9e-006                     vth0=0.42462821 k2=-0.0036779275              cit=0.00083837687              voff=-0.17771724 eta0=0.19777778                 etab=-0.034444444               u0=0.019857143 ua=-1.6811312e-009            ub=2.188862e-018              uc=8.0798373e-011 vsat=99665.553                  a0=1.4576238                  ags=2.3362286 keta=-0.056688151               pclm=0.68752834                 pdiblc2=0.0048541029 agidl=5.5747575e-011             tvoff=0.00101335                 kt1=-0.25720893 kt2=-0.03                      ute=-1.1959184                 ua1=1.5820317e-009 ub1=-1.8023129e-018            uc1=-5.1455782e-011            at=26962.815 lvth0=1.4681734e-010             lk2=7.7039341e-010             lcit=1.3669969e-010 lvoff=4.8102244e-009             lua=6.2492687e-017             lub=5.735946e-026 luc=3.4286804e-018             lvsat=-0.00078942563             la0=-4.3893092e-007 lags=-7.6142036e-008            lketa=8.4814293e-010             lpclm=-3.8469388e-008 lpdiblc2=-5.4833644e-010            lagidl=3.2223791e-017             ltvoff=2.05697e-010 lkt1=4.2163475e-009             lua1=-1.6163183e-016            lub1=7.2835374e-026 luc1=5.3344218e-018             lat=0.00029271504              lute=-1.0258503e-008 lu0=1.6157143e-009             wvth0=-5.638202e-009             wk2=-4.6394984e-009 wcit=5.8689796e-011             wvoff=-7.8583354e-009            weta0=-1.6e-007 wetab=-5e-009                    wua=-6.9165066e-017            wub=1.3198342e-025 wuc=5.1942347e-018             wa0=1.1672712e-006             wags=-5.2809826e-007 wketa=-2.4677684e-009            wpclm=1.122449e-008              wpdiblc2=-5.5824941e-009 wagidl=5.6023357e-017             wtvoff=1.70418e-011               wkt1=7.8453061e-009 wua1=-3.1589958e-016            wub1=2.2285714e-025             wuc1=1.4938776e-017 pvth0=1.3541588e-015             pk2=-3.1623067e-016            pcit=1.611098e-017 pvoff=-3.3819492e-015            pua=1.8407706e-023             pub=-6.4087596e-032 puc=-6.553164e-024             pa0=-2.7698391e-013            pags=6.2074247e-014 pketa=1.1850514e-015             ppclm=3.4622449e-014             ppdiblc2=2.0198854e-015 pagidl=-1.8889119e-023            ptvoff=-1.04848e-016              pkt1=1.6429506e-015 pua1=1.9586096e-022             pub1=-3.2314286e-032            puc1=3.9238775e-024 wat=-0.016082843               pat=1.7676944e-009             wvsat=0.0016922029 pvsat=-5.3408509e-010            wute=-3.6734694e-008            pute=9.2326531e-014 wu0=0                          pu0=0                          u0_mc=-2.22223e-05 vsat_mc=-131.519                   lvsat_mc=5.12925e-05                lu0_mc=-1.7e-18 wvsat_mc=0.00118367                 pvsat_mc=-4.61633e-10               wu0_mc=2e-10 pu0_mc=-3.5e-23 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.12 nmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=9e-007                     wmax=9e-006                     vth0=0.38425928 k2=0.0047360642               cit=0.00016771927              voff=-0.16697409 eta0=0.19777778                 etab=-0.034444444               u0=0.033866941 ua=-9.5360868e-010            ub=1.7989026e-018             uc=2.2002517e-010 vsat=96449.982                  a0=6.3598755                  ags=3.9039781 keta=-0.16123048                pclm=1.0672839                  pdiblc2=0.0061332682 agidl=9.6943678e-010             tvoff=0.00273223                 kt1=-0.24585524 kt2=-0.055369561               ute=-2.9868313                 ua1=-5.2226012e-010 ub1=-3.7368999e-018            uc1=-2.3714129e-010            at=19207.072 lvth0=6.0003127e-009             lk2=-4.4963537e-010            lcit=2.3394504e-010 lvoff=3.2524675e-009             lua=-4.2998077e-017            lub=1.1390357e-025 luc=-1.6759205e-017            lvsat=-0.0003231678              la0=-1.1497574e-006 lags=-3.0346571e-007            lketa=1.600678e-008              lpclm=-9.3533951e-008 lpdiblc2=-7.3381541e-010            lagidl=-1.0026114e-016            ltvoff=-4.35401e-011 lkt1=2.5700635e-009             lua1=1.4349048e-016             lub1=3.5335048e-025 luc1=3.225882e-017              lat=0.0014172976               lute=2.4942387e-007 lu0=-4.1570645e-010            lkt2=3.6785863e-009             wvth0=-1.2792961e-008 wk2=-2.8985751e-008            wcit=-1.565029e-009             wvoff=-1.5035255e-008 weta0=-1.6e-007                  wetab=-5e-009                    wua=-1.4765777e-015 wub=-2.0679012e-025            wuc=-1.601621e-016             wa0=4.9965424e-007 wags=-3.5802469e-007            wketa=6.557983e-008              wpclm=-2.1444444e-007 wpdiblc2=-2.5588303e-008            wagidl=-2.6582055e-016            wtvoff=-1.63204e-009 wkt1=3.4254963e-008             wua1=2.5401382e-015             wub1=1.4965432e-024 wuc1=1.4004938e-016             pvth0=2.3915988e-015             pk2=3.213976e-015 pcit=2.5155021e-016             pvoff=-2.3412958e-015            pua=2.2248254e-022 pub=-1.4965432e-032            puc=1.7423504e-023             pa0=-1.8017945e-013 pags=3.741358e-014              pketa=-8.6818503e-015            ppclm=6.7344444e-014 ppdiblc2=4.9207276e-015             pagidl=2.7778248e-023             ptvoff=1.34268e-016 pkt1=-2.1864496e-015            pua1=-2.1826452e-022            pub1=-2.1699876e-031 puc1=-1.4217161e-023            wat=-0.013223005               pat=1.353018e-009 wvsat=-0.0050028647              pvsat=4.3669973e-010             wute=2.1481481e-006 pute=-2.2448148e-013            wu0=-2.5802469e-008            pu0=3.741358e-015 wkt2=-3.8961728e-009            pkt2=5.6494506e-016             voff_mc=-0.00573388 u0_mc=-0.0001369                 vsat_mc=795.61                     lvoff_mc=8.31413e-10 lvsat_mc=-8.31413e-05               lu0_mc=1.66283e-11                wvoff_mc=5.16049e-09 pvoff_mc=-7.48272e-16               wvsat_mc=-0.00716049                pvsat_mc=7.48272e-10 wu0_mc=1.2321e-09                 pu0_mc=-1.49654e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.13 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=5.4e-007                   wmax=9e-007                     vth0=0.44265375 k2=0.015628011                cit=0.0002773125               voff=-0.19156542 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.477435e-009             ub=2.4e-018                   uc=9.945e-011 vsat=100000                     a0=2.0975732                  ags=0.75891614 keta=-0.060655368               pclm=0.2625                     pdiblc2=0.001025238 agidl=3.6634794e-010             tvoff=0.000855116                kt1=-0.19975742 kt2=-0.03                      ute=-1                         ua1=1.845236e-009 ub1=-1.425e-018                uc1=-2.375e-012                at=120000 lvth0=0                          lk2=0                          luc=0 lketa=0                          lpdiblc2=0                          lu0=0 wvth0=-8.434125e-009             wk2=-3.7770834e-009            wcit=8.0645625e-010 wvoff=1.4882778e-008             weta0=1.755e-007                 wetab=7.7274e-009 wua=-6.3659722e-017            wub=5.4e-026                   wuc=-6.075e-018 wa0=1.3104855e-009             wags=8.1996584e-009             wketa=5.3878817e-009 wpclm=-3.375e-008                wpdiblc2=-4.7142e-012               wagidl=4.3497655e-017 wtvoff=6.58876e-010               wkt1=-1.168722e-009             wua1=2.6330762e-016 wub1=-4.725e-025                wuc1=-1.92375e-017              pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.14 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=0.44529752 k2=0.016742369                cit=0.00012968253              voff=-0.1948109 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.4690192e-009            ub=2.3947771e-018             uc=9.9373205e-011 vsat=100275.25                  a0=2.1756294                  ags=0.67913341 keta=-0.055751144               pclm=0.26077967                 pdiblc2=0.00078132821 agidl=3.8013043e-010             tvoff=0.000736711                kt1=-0.19432055 kt2=-0.03                      ute=-1                         ua1=1.8143026e-009 ub1=-1.304577e-018             uc1=4.5235164e-012             at=119088.91 lvth0=-2.3820333e-008            lk2=-1.0040366e-008            lcit=1.330146e-009 lvoff=2.9241755e-008             lua=-7.5825805e-017            lub=4.7058479e-026 luc=6.9192705e-019             lvsat=-0.0024800252              la0=-7.0328661e-007 lags=7.1884237e-007             lketa=-4.4187057e-008            lpclm=1.5500158e-008 lpdiblc2=2.1976273e-009             lagidl=-1.2418024e-016            ltvoff=1.06683e-009 lkt1=-4.8986178e-008            lua1=2.7871022e-016             lub1=-1.085011e-024 luc1=-6.2155633e-017            lat=0.0082088836               lu0=0 wvth0=-9.0976935e-009            wk2=-3.775463e-009             wcit=9.3602536e-010 wvoff=1.7271149e-008             weta0=1.755e-007                 wetab=7.7274e-009 wua=-6.7425822e-017            wub=6.0536284e-026             wuc=-5.4262023e-018 wa0=-7.3966958e-009            wags=2.2535422e-008             wketa=3.5415951e-009 wpclm=-6.6264205e-008            wpdiblc2=1.6538302e-010             wagidl=5.8273177e-017 wtvoff=7.83165e-010               wkt1=-1.8327029e-009            wua1=3.3298884e-016 wub1=-5.9326705e-025            wuc1=-2.4672017e-017            pvth0=5.9787519e-015 pk2=-1.4599933e-017            pcit=-1.1674176e-015            pvoff=-2.1519221e-014 pua=3.393256e-023              pub=-5.889192e-032             puc=-5.8456675e-024 pa0=7.8451704e-014             pags=-1.2916523e-013            pketa=1.6635042e-014 ppclm=2.9295298e-013             ppdiblc2=-1.532576e-015             pagidl=-1.3312746e-022 ptvoff=-1.11984e-015              pkt1=5.9824682e-015             pua1=-6.2782784e-022 pub1=1.0881111e-030             puc1=4.8964999e-023             wat=0.0021329318 pat=-1.9217716e-008            wvsat=0                          wu0=0 pu0=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.15 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=0.41687939 k2=0.015027069                cit=0.0014922222               voff=-0.14124298 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.6691786e-009            ub=2.5914789e-018             uc=1.1317493e-010 vsat=98000                      a0=2.6758876                  ags=1.3561141 keta=-0.13521583                pclm=-0.57833333                pdiblc2=0.0071245349 agidl=4.6390646e-010             tvoff=0.00266137                 kt1=-0.25058004 kt2=-0.03                      ute=-1                         ua1=2.3680978e-009 ub1=-2.8333333e-018            uc1=-8.45e-011                 at=268625.78 lvth0=7.1554227e-009             lk2=-8.1706889e-009            lcit=-1.5502222e-010 lvoff=-2.9147278e-008            lua=1.4234791e-016             lub=-1.6734649e-025 luc=-1.4351957e-017            la0=-1.2485681e-006            lags=-1.9066563e-008 lketa=4.2429448e-008             lpclm=9.3013333e-007             lpdiblc2=-4.716468e-009 lagidl=-2.154961e-016             ltvoff=-1.03105e-009              lkt1=1.2336668e-008 lua1=-3.2492658e-016            lub1=5.8133333e-025             luc1=3.488e-017 lat=-0.1547863                 lu0=0                          wvth0=-2.2795517e-009 wk2=-2.1966346e-009            wcit=-1.35e-010                 wvoff=-8.9983344e-009 weta0=1.755e-007                 wetab=7.7274e-009                wua=5.5086963e-017 wub=-6.10386e-026              wuc=-1.196424e-017             wa0=-5.1557932e-007 wags=-3.2675515e-007            wketa=4.1481528e-008             wpclm=5.865e-007 wpdiblc2=-4.7292488e-009            wagidl=-1.4237869e-016            wtvoff=-6.43191e-010 wkt1=9.74604e-009               wua1=-3.32088e-016              wub1=6.93e-025 wuc1=4.137e-017                 pvth0=-1.4530227e-015            pk2=-1.7355228e-015 pcit=-1.8994406e-030            pvoff=7.1145155e-015             pua=-9.9606377e-023 pub=7.3624704e-032             puc=1.2807936e-024             pa0=6.3237077e-013 pags=2.5156149e-013             pketa=-2.4719484e-014            ppclm=-4.1856e-013 ppdiblc2=3.8025727e-015             pagidl=8.5583078e-023             ptvoff=4.34884e-016 pkt1=-6.6383616e-015            pua1=9.710592e-023              pub1=-3.1392e-031 puc1=-2.30208e-023              wat=-0.0541608                 pat=4.2142452e-008 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.16 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.42823758 k2=0.0074162525               cit=0.000704                   voff=-0.18830252 eta0=-0.175                     etab=-0.048586                  u0=0.024 ua=-1.3845577e-009            ub=2.3768e-018                uc=8.6293031e-011 vsat=98000                      a0=0.335                      ags=0.82358353 keta=-0.076892699               pclm=1.148                      pdiblc2=-0.0053070628 agidl=3.7786914e-011             tvoff=0.000364301                kt1=-0.23801824 kt2=-0.03                      ute=-1                         ua1=2.6341272e-009 ub1=-2.627e-018                uc1=-5.652e-011                at=48359.117 lvth0=-1.138176e-010             lk2=-3.2997666e-009            lcit=3.4944e-010 lvoff=9.7083018e-010             lua=-3.9809478e-017            lub=-2.9952e-026 luc=2.85246e-018               la0=2.496e-007                 lags=3.2175299e-007 lketa=5.1026455e-009             lpclm=-1.7472e-007               lpdiblc2=3.2397545e-009 lagidl=5.7220404e-017             ltvoff=4.39071e-010               lkt1=4.2971136e-009 lua1=-4.9518543e-016            lub1=4.4928e-025                luc1=1.69728e-017 lat=-0.013815635               lu0=0                          wvth0=-4.139516e-009 wk2=-3.1392832e-009            wcit=7.56e-011                  wvoff=2.5255733e-009 weta0=1.755e-007                 wetab=7.7274e-009                wua=-1.750348e-016 wub=1.3824e-025                wuc=-1.7555231e-018            wa0=1.39914e-006 wags=5.3957483e-008             wketa=-6.6266894e-009            wpclm=-1.728e-007 wpdiblc2=3.1034139e-009             wagidl=3.0773946e-017             wtvoff=4.14658e-010 wkt1=6.820416e-009              wua1=-4.7601292e-016            wub1=4.9734e-025 wuc1=9.612e-018                 pvth0=-2.6264549e-016            pk2=-1.1322277e-015 pcit=-1.34784e-016              pvoff=-2.6078548e-016            pua=4.7671551e-023 pub=-5.39136e-032              puc=-5.2527852e-024            pa0=-5.930496e-013 pags=7.9054051e-015             pketa=6.0697748e-015             ppclm=6.7392e-014 ppdiblc2=-1.2103314e-015            pagidl=-2.5234608e-023            ptvoff=-2.42139e-016 pkt1=-4.7659622e-015            pua1=1.8921787e-022             pub1=-1.886976e-031 puc1=-2.69568e-024              wat=0.027186966                pat=-9.9201184e-009 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0                          u0_mc=-0.000312 lu0_mc=1.9968e-10                 wu0_mc=0.0                        pu0_mc=0.0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.17 nmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.4278394 k2=0.0016137502               cit=0.00087529592              voff=-0.1893543 eta0=-0.175                     etab=-0.048586                  u0=0.019857143 ua=-1.7426736e-009            ub=2.4242857e-018             uc=1.1704793e-010 vsat=106164.86                  a0=3.8942246                  ags=0.99673701 keta=-0.075270054               pclm=0.54020408                 pdiblc2=-0.0080268894 agidl=1.9167852e-010             tvoff=0.00132648                 kt1=-0.24353592 kt2=-0.03                      ute=-1.5918367                 ua1=4.6462701e-010 ub1=-1.3122449e-018            uc1=-6.0938775e-011            at=7534.9734 lvth0=4.1472154e-011             lk2=-1.0367907e-009            lcit=2.8263459e-010 lvoff=1.3810247e-009             lua=9.9855737e-017             lub=-4.8471429e-026 luc=-9.1419495e-018            lvsat=-0.003184294               la0=-1.1384976e-006 lags=2.5422313e-007             lketa=4.4698141e-009             lpclm=6.2320408e-008 lpdiblc2=4.3004868e-009             lagidl=-2.7973237e-018            ltvoff=6.38207e-011 lkt1=6.4490082e-009             lua1=3.5091965e-016             lub1=-6.347449e-026 luc1=1.8696122e-017             lat=0.0021057812               lute=2.3081633e-007 lu0=1.6157143e-009             wvth0=-8.5282722e-009            wk2=-9.4020082e-009 wcit=2.5462653e-011             wvoff=2.6150196e-009             weta0=1.755e-007 wetab=7.7274e-009                wua=-1.3776875e-017            wub=-7.9897959e-026 wuc=-2.7430364e-017            wa0=-1.0256695e-006            wags=6.7744418e-007 wketa=1.4255945e-008             wpclm=1.4381633e-007             wpdiblc2=6.0103989e-009 wagidl=-6.6314496e-017            wtvoff=-2.64778e-010              wkt1=-4.4604e-009 wua1=6.8976465e-016             wub1=-2.1820408e-025            wuc1=2.3473469e-017 pvth0=1.4489694e-015             pk2=1.310235e-015              pcit=-1.1523044e-016 pvoff=-2.9566952e-016            pua=-1.5219039e-023            pub=3.1160204e-032 puc=4.7604028e-024             pa0=3.5262611e-013             pags=-2.3525441e-013 pketa=-2.0744527e-015            ppclm=-5.6088367e-014            ppdiblc2=-2.3440556e-015 pagidl=1.2629884e-023             ptvoff=2.28404e-017               pkt1=-3.66444e-016 pua1=-2.6543538e-022            pub1=9.0364592e-032             puc1=-8.1016531e-024 wat=0.0014022142               pat=1.359349e-010              wvsat=-0.0041571703 pvsat=1.6212964e-009             wute=3.1959184e-007             pute=-1.2464082e-013 wu0=0                          pu0=0                          u0_mc=2.2449e-05 vsat_mc=1627.55                    lvsat_mc=-0.000634743               lu0_mc=6.92451e-11 wvsat_mc=-0.000399491               pvsat_mc=1.55801e-10                wu0_mc=1.59796e-10 pu0_mc=-6.23204e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.18 nmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.3410019 k2=-0.020073327               cit=-0.00069857043             voff=-0.16658705 eta0=-0.36851852                etab=-0.048586659               u0=-0.041246914 ua=-5.2215322e-009            ub=1.4191358e-018             uc=-4.966142e-011 vsat=62228.783                  a0=4.8774446                  ags=7.2654321 keta=-0.091336901               pclm=1.0174159                  pdiblc2=-0.032213879 agidl=5.9138425e-010             tvoff=0.00161713                 kt1=-0.19038521 kt2=-0.065542901               ute=1.5481482                  ua1=5.3059996e-009 ub1=-2.407963e-018             uc1=-3.0049383e-011            at=2114.167 lvth0=1.263291e-008              lk2=2.1078354e-009             lcit=5.1084521e-010 lvoff=-1.9202269e-009            lua=6.0429024e-016             lub=9.7275309e-026 luc=1.5030906e-017             lvsat=0.0031864367               la0=-1.2810645e-006 lags=-6.5473765e-007            lketa=6.7995069e-009             lpclm=-6.8753056e-009 lpdiblc2=7.8076004e-009             lagidl=-6.0754654e-017            ltvoff=2.16765e-011 lkt1=-1.2578446e-009            lua1=-3.5107937e-016            lub1=9.540463e-026 luc1=1.4217161e-017             lat=0.0028917981               lute=-2.2448148e-007 lu0=1.0475803e-008             lkt2=5.1537207e-009             wvth0=2.6138683e-008 wk2=-6.6572997e-009            wcit=-7.8536828e-010            wvoff=-1.5383592e-008 weta0=3.4966667e-007             wetab=7.7279932e-009             wua=2.3645535e-015 wub=1.35e-025                  wuc=8.2555833e-017             wa0=1.8338421e-006 wags=-3.3833333e-006            wketa=2.6756132e-009             wpclm=-1.695632e-007 wpdiblc2=8.9241302e-009             wagidl=7.4426721e-017             wtvoff=-6.28451e-010 wkt1=-1.5668067e-008            wua1=-2.7052955e-015            wub1=3.005e-025 wuc1=-4.6333333e-017            pvth0=-3.5777391e-015            pk2=9.1225229e-016 pcit=2.3400511e-018             pvoff=2.3141292e-015             pua=-3.6007694e-022 pub=3.9305792e-045             puc=-1.1187596e-023            pa0=-6.200307e-014 pags=3.5355833e-013             pketa=-3.9530453e-016            ppclm=-1.0648336e-014 ppdiblc2=-2.7665466e-015            pagidl=-7.7775924e-024            ptvoff=7.55731e-017 pkt1=1.2586677e-015             pua1=2.2684835e-022             pub1=1.51525e-032 puc1=2.0203333e-024             wat=0.0021606097               pat=2.5967546e-011 wvsat=0.025796214                pvsat=-2.7219443e-009            wute=-1.9333333e-006 pute=2.0203333e-013             wu0=4.18e-008                  pu0=-6.061e-015 wkt2=5.2598333e-009             pkt2=-7.6267583e-016            leta0=2.8060185e-008 peta0=-2.5254167e-014            letab=9.5572991e-014             petab=-8.6015692e-020 u0_mc=0.00308024                 vsat_mc=-17586.4                   lvsat_mc=0.00215128 lu0_mc=-3.74136e-10               wvsat_mc=0.00938334                 pvsat_mc=-1.26271e-09 wu0_mc=-1.66333e-09               pu0_mc=2.02034e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.19 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.42910039 k2=0.016243241                cit=0.00135265                 voff=-0.1681236 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.6175468e-009            ub=2.62e-018                  uc=1.0786e-010 vsat=100000                     a0=2.3                        ags=0.87190207 keta=-0.07279409                pclm=0.2                        pdiblc2=0.001133524 agidl=6.4044621e-010             tvoff=0.00209897                 kt1=-0.20486516 kt2=-0.03                      ute=-1                         ua1=2.764928e-009 ub1=-2.9e-018                  uc1=-5.8e-011                  at=120000 lvth0=0                          lk2=0                          luc=0 lketa=0                          lpdiblc2=0                          lu0=0 wvth0=-1.1153117e-009            wk2=-4.1093078e-009            wcit=2.25774e-010 wvoff=2.2241952e-009             weta0=-8.64e-008                 wetab=1.001808e-008 wua=1.200069e-017              wub=-6.48e-026                 wuc=-1.06164e-017 wa0=-1.08e-007                 wags=-5.2812744e-008            wketa=1.1942791e-008 wpdiblc2=-6.318864e-011             wagidl=-1.0451541e-016            wtvoff=-1.28045e-011 wkt1=1.5894576e-009             wua1=-2.3332609e-016            wub1=3.24e-025 wuc1=1.08e-017                  pvth0=0                          pk2=0 puc=0                          pketa=0                          wvsat=0 wu0=0                          pu0=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.20 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.43046267 k2=0.016946903                cit=0.001359896                voff=-0.16659847 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.6215494e-009            ub=2.6441204e-018             uc=1.0860848e-010 vsat=100275.25                  a0=2.3756944                  ags=0.85336935 keta=-0.073629861               pclm=0.16240051                 pdiblc2=0.0011381378 agidl=7.2765024e-010             tvoff=0.00224871                 kt1=-0.19934563 kt2=-0.03                      ute=-1                         ua1=2.9306917e-009 ub1=-3.1050631e-018            uc1=-6.4479444e-011            at=124475.61 lvth0=-1.2274131e-008            lk2=-6.3399888e-009            lcit=-6.5286665e-011 lvoff=-1.3741403e-008            lua=3.6062828e-017             lub=-2.1732461e-025 luc=-6.7438087e-018            lvsat=-0.0024800252              la0=-6.8200694e-007 lags=1.6697981e-007             lketa=7.5302965e-009             lpclm=3.3877145e-007 lpdiblc2=-4.1570183e-011            lagidl=-7.8570829e-016            ltvoff=-1.34919e-009 lkt1=-4.9731004e-008            lua1=-1.4935308e-015            lub1=1.8476188e-024 luc1=5.8379794e-017             lat=-0.040325211               lu0=0 wvth0=-1.0868769e-009            wk2=-3.8859112e-009            wcit=2.7171007e-010 wvoff=2.0364389e-009             weta0=-8.64e-008                 wetab=1.001808e-008 wua=1.4940457e-017             wub=-7.4109096e-026            wuc=-1.0413251e-017 wa0=-1.1543182e-007            wags=-7.1551984e-008            wketa=1.3196102e-008 wpclm=-1.3139454e-008            wpdiblc2=-2.7294147e-011            wagidl=-1.2938752e-016 wtvoff=-3.33155e-011              wkt1=8.8083671e-010             wua1=-2.6986131e-016 wub1=3.7899545e-025             wuc1=1.2589582e-017             pvth0=-2.5619692e-016 pk2=-2.0128038e-015            pcit=-4.1388397e-016            pvoff=1.6916839e-015 pua=-2.6487302e-023            pub=8.387495e-032              puc=-1.8303702e-024 pa0=6.6960682e-014             pags=1.6884055e-013             pketa=-1.1292329e-014 ppclm=1.1838649e-013             ppdiblc2=-3.2340938e-016            pagidl=2.2409769e-022 ptvoff=1.84804e-016               pkt1=6.3846742e-015             pua1=3.291823e-022 pub1=-4.9550905e-031            puc1=-1.6124132e-023            wat=-0.00077588182 pat=6.9906952e-009             wvsat=0                          wu0=0 pu0=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.21 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.40825089 k2=0.026188636                cit=0.0023170222               voff=-0.14985865 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.5635028e-009            ub=2.3803702e-018             uc=1.2319627e-010 vsat=98000                      a0=1.9633333                  ags=0.22111143 keta=-0.057600561               pclm=0.50619556                 pdiblc2=-0.00018 agidl=-2.0011244e-010            tvoff=0.00155439                 kt1=-0.26821861 kt2=-0.03                      ute=-1                         ua1=1.5935893e-009 ub1=-1.0686667e-018            uc1=5.4688666e-012             at=121763.2 lvth0=1.1936711e-008             lk2=-1.6413478e-008            lcit=-1.1085542e-009 lvoff=-3.1987806e-008            lua=-2.7207919e-017            lub=7.0163058e-026 luc=-2.2644499e-017            la0=-2.3253333e-007            lags=8.5614093e-007 lketa=-9.9416399e-009            lpclm=-3.5965156e-008            lpdiblc2=1.3952e-009 lagidl=2.2555302e-016             ltvoff=-5.92375e-010              lkt1=2.5340552e-008 lua1=-3.6089173e-017            lub1=-3.7205333e-025            luc1=-1.7863865e-017 lat=-0.037368688               lu0=0                          wvth0=2.37984e-009 wk2=-8.2238811e-009            wcit=-5.8039199e-010            wvoff=-4.3458699e-009 weta0=-8.64e-008                 wetab=1.001808e-008              wua=-1.9779576e-018 wub=5.296008e-026              wuc=-1.7375762e-017            wa0=-1.308e-007 wags=2.8614629e-007             wketa=-4.307161e-010             wpclm=8.544e-010 wpdiblc2=-7.848e-010                wagidl=2.1619151e-016             wtvoff=-4.54198e-011 wkt1=1.9270867e-008             wua1=8.614656e-017              wub1=-2.5992e-025 wuc1=-7.2131879e-018            pvth0=-4.0349184e-015            pk2=2.7155834e-015 pcit=5.1490727e-016             pvoff=8.6484006e-015             pua=-8.04623e-024 pub=-5.4630451e-032            puc=5.7587661e-024             pa0=8.3712e-014 pags=-2.2105056e-013            pketa=3.5609032e-015             ppclm=1.0313318e-013 ppdiblc2=5.02272e-016               pagidl=-1.5258345e-022            ptvoff=1.97998e-016 pkt1=-1.3660459e-014            pua1=-5.8866278e-023            pub1=2.009088e-031 puc1=5.4608869e-024             wat=0.025144992                pat=-2.1263057e-008 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0                          u0_mc=0.000284444 lu0_mc=-3.10044e-10               wu0_mc=-1.536e-10                 pu0_mc=1.67424e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.22 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.42382441 k2=0.011945321                cit=-3.7094974e-005            voff=-0.20219733 eta0=0.31                       etab=-0.052828                  u0=0.024 ua=-1.6241451e-009            ub=2.6928e-018                uc=1.0987428e-010 vsat=98000                      a0=2.146                      ags=2.0811878 keta=-0.09597384                pclm=0.4032                     pdiblc2=-0.00268 agidl=3.2981508e-010             tvoff=0.000731214                kt1=-0.21719232 kt2=-0.03                      ute=-1                         ua1=2.0848255e-009 ub1=-2.43e-018                 uc1=-6.993516e-011             at=142692.69 lvth0=1.9696595e-009             lk2=-7.2977563e-009            lcit=3.9808079e-010 lvoff=1.5089478e-009             lua=1.1603155e-017             lub=-1.29792e-025 luc=-1.4118427e-017            la0=-3.4944e-007               lags=-3.3430793e-007 lketa=1.4617258e-008             lpclm=2.9952e-008                lpdiblc2=2.9952e-009 lagidl=-1.1360058e-016            ltvoff=-6.5545e-011               lkt1=-7.3162752e-009 lua1=-3.5048033e-016            lub1=4.992e-025                 luc1=3.0394712e-017 lat=-0.050763563               lu0=0                          wvth0=-1.7564026e-009 wk2=-5.5849801e-009            wcit=4.7579129e-010             wvoff=1.002877e-008 weta0=-8.64e-008                 wetab=1.001808e-008              wua=-4.5657581e-017 wub=-3.24e-026                 wuc=-1.4489399e-017            wa0=4.212e-007 wags=-6.2514881e-007            wketa=3.6771267e-009             wpclm=2.29392e-007 wpdiblc2=1.6848e-009                wagidl=-1.2692126e-016            wtvoff=2.16525e-010 wkt1=-4.4255808e-009            wua1=-1.7938999e-016            wub1=3.9096e-025 wuc1=1.6856186e-017             pvth0=-1.3877231e-015            pk2=1.0266867e-015 pcit=-1.6105003e-016            pvoff=-5.51369e-016              pua=1.9908729e-023 pub=-1.7913775e-045            puc=3.9114937e-024             pa0=-2.69568e-013 pags=3.621783e-013              pketa=9.3188385e-016             ppclm=-4.313088e-014 ppdiblc2=-1.078272e-015             pagidl=6.7008726e-023             ptvoff=3.03534e-017 pkt1=1.5052677e-015             pua1=1.1107711e-022             pub1=-2.156544e-031 puc1=-9.9435127e-024            wat=-0.023753164               pat=1.0031763e-008 wvsat=0                          wu0=0                          pu0=0 pvsat=0                          lvsat=0                          u0_mc=-0.000824 lu0_mc=3.9936e-10                 wu0_mc=2.7648e-10                 pu0_mc=-1.07827e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.23 nmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.42673106 k2=-0.0093237196              cit=0.001092301                voff=-0.20711602 eta0=0.31                       etab=-0.052828                  u0=0.019857143 ua=-1.641151e-009             ub=2.1469388e-018             uc=6.8745074e-011 vsat=98200.608                  a0=1.8721589                  ags=1.8300216 keta=-0.073219292               pclm=0.66938775                 pdiblc2=0.010515236 agidl=-5.3456526e-011            tvoff=0.000157831                kt1=-0.24776033 kt2=-0.03                      ute=-0.52653061                ua1=2.5336766e-009 ub1=-1.7122449e-018            uc1=2.6086531e-011             at=2788.9622 lvth0=8.3606567e-010             lk2=9.971694e-010              lcit=-4.2383648e-011 lvoff=3.4272386e-009             lua=1.8235438e-017             lub=8.3093878e-026 luc=1.9219643e-018             lvsat=-7.823704e-005             la0=-2.4264198e-007 lags=-2.3635314e-007            lketa=5.7429849e-009             lpclm=-7.3861224e-008 lpdiblc2=-2.1509422e-009            lagidl=3.5875339e-017             ltvoff=1.58075e-010 lkt1=4.6052474e-009             lua1=-5.2553226e-016            lub1=2.1927551e-025 luc1=-7.0537469e-018            lat=0.0037988918               lute=-1.8465306e-007 lu0=1.6157143e-009             wvth0=-7.9297669e-009            wk2=-3.4957746e-009 wcit=-9.1720102e-011            wvoff=1.220635e-008              weta0=-8.64e-008 wetab=1.001808e-008              wua=-6.8599102e-017            wub=6.9869388e-026 wuc=-1.3468234e-018            wa0=6.6245972e-008             wags=2.2747047e-007 wketa=1.3148534e-008             wpclm=7.4057143e-008             wpdiblc2=-4.002349e-009 wagidl=6.605843e-017              wtvoff=3.66294e-010               wkt1=-2.1792196e-009 wua1=-4.2752214e-016            wub1=-2.2040816e-027            wuc1=-2.3520196e-017 pvth0=1.0198889e-015             pk2=2.1189658e-016             pcit=6.0279415e-017 pvoff=-1.400625e-015             pua=2.8855922e-023             pub=-3.9885061e-032 puc=-1.2141106e-024            pa0=-1.3113593e-013            pags=2.9656782e-014 pketa=-2.7619649e-015            ppclm=1.7449714e-014             ppdiblc2=1.1397161e-015 pagidl=-8.2533537e-024            ptvoff=-2.80566e-017              pkt1=6.2918684e-016 pua1=2.0784865e-022             pub1=-6.2320408e-032            puc1=5.8032764e-024 wat=0.0039650602               pat=-7.783448e-010             wvsat=0.0001435239 pvsat=-5.5974321e-011            wute=-2.5567347e-007            pute=9.9712653e-014 wu0=0                          pu0=0                          u0_mc=0.000318367 vsat_mc=2071.43                    lvsat_mc=-0.000807854               lu0_mc=-4.61635e-11 wvsat_mc=-0.000639184               pvsat_mc=2.49281e-10                wu0_mc=-2.7e-16 pu0_mc=-2.7e-23 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.24 nmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=0.40648154 k2=-0.028089147               cit=-0.0071268385              voff=-0.23427534 eta0=0.85185185                 etab=-0.052826682               u0=0.046481482 ua=7.8899628e-010             ub=5.0098765e-019             uc=1.0518916e-010 vsat=123371.75                  a0=15.70361                   ags=-2.3802469 keta=-0.089616651               pclm=-0.16189353                pdiblc2=-0.025783529 agidl=6.6862081e-010             tvoff=-0.0012084                 kt1=-0.20785674 kt2=-0.055802469               ute=-4.8962963                 ua1=-4.3428677e-009 ub1=-2.7544444e-018            uc1=-3.078321e-010             at=7717.1282 lvth0=3.7722463e-009             lk2=3.7181564e-009             lcit=1.1493916e-009 lvoff=7.3653392e-009             lua=-3.3413591e-016            lub=3.2175679e-025 luc=-3.3624286e-018            lvsat=-0.0037280531              la0=-2.2482024e-006 lags=3.741358e-007              lketa=8.1206019e-009             lpclm=4.6674562e-008 lpdiblc2=3.1123788e-009             lagidl=-6.8825874e-017            ltvoff=3.56177e-010 lkt1=-1.1807726e-009            lua1=4.7156667e-016             lub1=3.7039444e-025 luc1=4.1364454e-017             lat=0.0030843077               lute=4.4896296e-007 lu0=-2.2448148e-009            lkt2=3.741358e-009              wvth0=-9.2203222e-009 wk2=-2.3287568e-009            wcit=2.6858965e-009             wvoff=2.1168084e-008 weta0=-3.0933333e-007            wetab=1.0017605e-008             wua=-8.811319e-016 wub=6.308e-025                 wuc=-1.0634811e-018            wa0=-4.0122871e-006 wags=1.8253333e-006             wketa=1.7466781e-009             wpclm=4.6726389e-007 wpdiblc2=5.4517409e-009             wagidl=3.2718979e-017             wtvoff=8.97333e-010 wkt1=-6.23344e-009              wua1=2.5050928e-015             wub1=4.876e-025 wuc1=1.0366933e-016             pvth0=1.2070195e-015             pk2=4.2679e-017 pcit=-3.4247499e-016            pvoff=-2.7000765e-015            pua=1.4667318e-022 pub=-1.2122e-031               puc=-1.2551952e-024            pa0=4.6025137e-013 pags=-2.0203333e-013            pketa=-1.1086958e-015            ppclm=-3.9565264e-014 ppdiblc2=-2.3112693e-016            pagidl=-3.4191333e-024            ptvoff=-1.05057e-016 pkt1=1.2170488e-015             pua1=-2.1738051e-022            pub1=-1.33342e-031 puc1=-1.2639205e-023            wat=-0.00086498939             pat=-7.7987614e-011 wvsat=-0.0072209897              pvsat=1.0118802e-009             wute=1.5466667e-006 pute=-1.6162667e-013            wu0=-5.5733333e-009            pu0=8.0813333e-016 leta0=-7.8568518e-008            peta0=3.2325333e-014             letab=-1.9114598e-013 petab=6.8812553e-020             vsat_mc=-2209.86                   lvsat_mc=-0.000187069 wvsat_mc=0.00108                    pvsat_mc=-6.7e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.25 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.39330752 k2=0.0076464838               cit=0.002299                   voff=-0.15436512 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-1.865698e-009             ub=2.4e-018                   uc=5.4471019e-011 vsat=100000                     a0=1.2                        ags=0.572 keta=-0.03187431                pclm=0.30304                    pdiblc2=0.000838 agidl=-5.41322e-013              tvoff=0.0023061                  kt1=-0.21177 kt2=-0.03                      ute=-1                         ua1=1.7432e-009 ub1=-1.68e-018                 uc1=-1.2e-011                  at=120000 lvth0=0                          lk2=0                          luc=0 lketa=0                          lpdiblc2=0                          lu0=0 wvth0=1.1770122e-008             wk2=-1.0144751e-009            wcit=-1.14912e-010 wvoff=-2.7288576e-009            weta0=1.152e-007                 wetab=1.4688e-008 wua=1.013351e-016              wub=1.44e-026                  wuc=8.6036332e-018 wa0=2.88e-007                  wags=5.5152e-008                wketa=-2.7883292e-009 wpclm=-3.70944e-008              wpdiblc2=4.32e-011                  wagidl=1.262401e-016 wtvoff=-8.7372e-011               wkt1=4.0752e-009                wua1=1.34496e-016 wub1=-1.152e-025                wuc1=-5.76e-018                 pvth0=0 pk2=0                          puc=0                          pketa=0 wvsat=0                          wu0=2.88e-009                  pu0=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.26 nmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.39272144 k2=0.0096380468               cit=0.0024777765               voff=-0.14973871 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-1.8291497e-009            ub=2.3637836e-018             uc=5.488193e-011 vsat=100275.25                  a0=1.0098155                  ags=0.54445742 keta=-0.0310503                 pclm=0.16693313                 pdiblc2=0.0013662096 agidl=-3.6673871e-011            tvoff=0.00259595                 kt1=-0.20323417 kt2=-0.03                      ute=-1                         ua1=1.8738701e-009 ub1=-1.842399e-018             uc1=-1.6789394e-011            at=116404.45 lvth0=5.280569e-009              lk2=-1.7943983e-008            lcit=-1.6107764e-009 lvoff=-4.1683917e-008            lua=-3.2929969e-016            lub=3.2630932e-025 luc=-3.7023136e-018            lvsat=-0.0024800252              la0=1.7135619e-006 lags=2.4815862e-007             lketa=-7.4243277e-009            lpclm=1.2263229e-006 lpdiblc2=-4.7591685e-009            lagidl=3.2555427e-016             ltvoff=-2.61158e-009 lkt1=-7.6907865e-008            lua1=-1.1773374e-015            lub1=1.4632149e-024 luc1=4.3152439e-017             lat=0.032395875                lu0=0 wvth0=1.2499966e-008             wk2=-1.2547231e-009            wcit=-1.3072691e-010 wvoff=-4.0330739e-009            weta0=1.152e-007                 wetab=1.4688e-008 wua=8.9676591e-017             wub=2.6812127e-026             wuc=8.9283068e-018 wa0=3.7628459e-007             wags=3.9656308e-008             wketa=-2.1325396e-009 wpclm=-1.47712e-008              wpdiblc2=-1.094e-010                wagidl=1.4576916e-016 wtvoff=-1.58323e-010              wkt1=2.2807112e-009             wua1=1.1059448e-016 wub1=-7.5563636e-026            wuc1=-4.5788364e-018            pvth0=-6.5758889e-015 pk2=2.1646339e-015             pcit=1.4249233e-016             pvoff=1.1750989e-014 pua=1.050432e-022              pub=-1.1183327e-031            puc=-2.9253085e-024 pa0=-7.9544412e-013            pags=1.3961618e-013             pketa=-5.908664e-015 ppclm=-2.0113203e-013            ppdiblc2=1.374926e-015              pagidl=-1.7595683e-022 ptvoff=6.39265e-016               pkt1=1.6168344e-014             pua1=2.153527e-022 pub1=-3.5712364e-031            puc1=-1.0642284e-023            wat=0.0021297332 pat=-1.9188896e-008            wvsat=0                          wu0=2.88e-009 pu0=0                          pvsat=0                          u0_mc=8.25758e-05 lu0_mc=-7.44008e-10               wu0_mc=-2.97273e-11               pu0_mc=2.67843e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.27 nmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.40147711 k2=-0.0019638134              cit=0.0025840223               voff=-0.17473404 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-2.3847245e-009            ub=3.0942967e-018             uc=5.3452918e-011 vsat=98000                      a0=3.4094686                  ags=1.3700218 keta=-0.097546714               pclm=1.0530667                  pdiblc2=-0.0035688889 agidl=7.4696333e-010             tvoff=0.000470243                kt1=-0.30130308 kt2=-0.03                      ute=-1                         ua1=8.9151324e-010 ub1=-7.8444444e-019            uc1=5.2227834e-011             at=307500.29 lvth0=-4.2631111e-009            lk2=-5.2979549e-009            lcit=-1.7265843e-009 lvoff=-1.4439018e-008            lua=2.7627682e-016             lub=-4.6994987e-025 luc=-2.1446897e-018            la0=-9.0205992e-007            lags=-6.5170654e-007 lketa=6.5056763e-008             lpclm=2.6043733e-007             lpdiblc2=6.2008889e-010 lagidl=-5.2861028e-016            ltvoff=-2.94555e-010              lkt1=2.9987251e-008 lua1=-1.0656848e-016            lub1=3.1004444e-025             luc1=-3.2076339e-017 lat=-0.17589858                lu0=0                          wvth0=4.8184e-009 wk2=1.9110007e-009             wcit=-6.7651201e-010            wvoff=4.6092676e-009 weta0=1.152e-007                 wetab=1.4688e-008                wua=2.9366186e-016 wub=-2.0405344e-025            wuc=7.7318451e-018             wa0=-6.5140871e-007 wags=-1.2746144e-007            wketa=1.3949899e-008             wpclm=-1.960192e-007 wpdiblc2=4.352e-010                 wagidl=-1.2475576e-016            wtvoff=3.44872e-010 wkt1=3.1181275e-008             wua1=3.3889395e-016             wub1=-3.6224e-025 wuc1=-2.4046416e-017            pvth0=1.7970176e-015             pk2=-1.286005e-015 pcit=7.3739809e-016             pvoff=2.3308367e-015             pua=-1.1730074e-022 pub=1.398102e-031              puc=-1.6211653e-024            pa0=3.2474157e-013 pags=3.2177453e-013             pketa=-2.3438522e-014            ppclm=-3.571712e-015 ppdiblc2=7.81312e-016               pagidl=1.1891534e-022             ptvoff=9.07828e-017 pkt1=-1.533327e-014             pua1=-3.3493729e-023            pub1=-4.46464e-032 puc1=1.0577377e-023             wat=-0.04172036                pat=2.8607705e-008 wvsat=0                          wu0=2.88e-009                  pu0=0 pvsat=0                          lvsat=0                          u0_mc=-0.00131111 lu0_mc=7.75107e-10                wu0_mc=4.208e-10                  pu0_mc=-2.23232e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.28 nmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.37668621 k2=-0.0088550293              cit=-0.0011503126              voff=-0.18279738 eta0=-0.25                      etab=-0.0658                    u0=0.016 ua=-2.2657003e-009            ub=2.75e-018                  uc=4.960161e-011 vsat=98000                      a0=4.652                      ags=2.1863257 keta=-0.013461155               pclm=1.4756                     pdiblc2=0.00055315936 agidl=-7.7738591e-010            tvoff=0.00048736                 kt1=-0.21043728 kt2=-0.03                      ute=-1                         ua1=1.9438707e-011 ub1=1.104e-018                 uc1=6.7797899e-011             at=44869.759 lvth0=1.1603065e-008             lk2=-8.875767e-010             lcit=6.6339003e-010 lvoff=-9.2784757e-009            lua=2.0010133e-016             lub=-2.496e-025 luc=3.2014694e-019             la0=-1.69728e-006              lags=-1.1741411e-006 lketa=1.1242006e-008             lpclm=-9.984e-009                lpdiblc2=-2.018022e-009 lagidl=4.4697323e-016             ltvoff=-3.0551e-010               lkt1=-2.8166861e-008 lua1=4.5155923e-016             lub1=-8.9856e-025               luc1=-4.2041181e-017 lat=-0.0078150459              lu0=0                          wvth0=1.5213348e-008 wk2=1.9031459e-009             wcit=8.7654962e-010             wvoff=3.0447884e-009 weta0=1.152e-007                 wetab=1.4688e-008                wua=1.8530229e-016 wub=-5.2992e-026               wuc=7.2087633e-018             wa0=-4.8096e-007 wags=-6.6299847e-007            wketa=-2.602744e-008             wpclm=-1.56672e-007 wpdiblc2=5.2086263e-010             wagidl=2.7167109e-016             wtvoff=3.04312e-010 wkt1=-6.8573952e-009            wua1=5.6414926e-016             wub1=-8.8128e-025 wuc1=-3.2727715e-017            pvth0=-4.8557492e-015            pk2=-1.2809779e-015 pcit=-2.5656135e-016            pvoff=3.3321034e-015             pua=-4.7950612e-023 pub=4.313088e-032              puc=-1.2863929e-024            pa0=2.156544e-013 pags=6.6451823e-013             pketa=2.1469748e-015             ppclm=-2.875392e-014 ppdiblc2=7.2648792e-016             pagidl=-1.3479785e-022            ptvoff=1.16741e-016 pkt1=9.0114785e-015             pua1=-1.7765713e-022            pub1=2.875392e-031 puc1=1.6133409e-023             wat=0.011463092                pat=-5.4297033e-009 wvsat=0                          wu0=2.88e-009                  pu0=0 pvsat=0                          lvsat=0                          u0_mc=-0.00088 lu0_mc=4.992e-10                  wu0_mc=2.9664e-10                 pu0_mc=-1.43769e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.29 nmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.38352036 k2=-0.010941318               cit=-0.00036625255             voff=-0.19906137 eta0=-0.25                      etab=-0.0658                    u0=0.007122449 ua=-1.9391147e-009            ub=1.6838776e-018             uc=3.5876633e-011 vsat=97708.279                  a0=2.5176122                  ags=-3.5611185 keta=0.020332674                pclm=1.6571429                  pdiblc2=-0.018474406 agidl=3.8673953e-010             tvoff=-0.000591918               kt1=-0.3122542 kt2=-0.03                      ute=-1.2367347                 ua1=3.9997129e-010 ub1=-6.0816327e-019            uc1=-7.5746939e-011            at=27976.71 lvth0=8.9377483e-009             lk2=-7.3924006e-011            lcit=3.5760662e-010 lvoff=-2.9355197e-009            lua=7.273293e-017              lub=1.6618776e-025 luc=5.6728883e-018             lvsat=0.00011377115              la0=-8.6486878e-007 lags=1.0673622e-006             lketa=-1.9375876e-009            lpclm=-8.0785714e-008 lpdiblc2=5.4027286e-009             lagidl=-7.0356858e-018            ltvoff=1.15408e-010 lkt1=1.154174e-008              lua1=3.0315152e-016             lub1=-2.3081633e-025 luc1=1.3941306e-017             lat=-0.0012267567              lute=9.2326531e-008 lu0=3.4622449e-009             wvth0=7.6260855e-009             wk2=-2.913439e-009 wcit=4.3335918e-010             wvoff=9.3066741e-009             weta0=1.152e-007 wetab=1.4688e-008                wua=3.8667833e-017             wub=2.3657143e-025 wuc=1.0485816e-017             wa0=-1.6611722e-007            wags=2.1682809e-006 wketa=-2.0530174e-008            wpclm=-2.8153469e-007            wpdiblc2=6.4339224e-009 wagidl=-9.2412149e-017            wtvoff=6.36204e-010               wkt1=2.1038576e-008 wua1=3.4061178e-016             wub1=-3.9967347e-025            wuc1=1.3139853e-017 pvth0=-1.8967168e-015            pk2=5.974902e-016              pcit=-8.3717082e-017 pvoff=8.89968e-016               pua=9.2368251e-024             pub=-6.9798857e-032 puc=-2.5644433e-024            pa0=9.2865718e-014             pags=-4.3968073e-013 pketa=3.0412359e-018             ppclm=1.9942531e-014             ppdiblc2=-1.5796054e-015 pagidl=7.1946152e-024             ptvoff=-1.26967e-017              pkt1=-1.8679504e-015 pua1=-9.047751e-023             pub1=9.9712653e-032             puc1=-1.7549427e-024 wat=-0.005102529               pat=1.0308886e-009             wvsat=0.00032076222 pvsat=-1.2509727e-010            wu0=4.5844898e-009             pu0=-6.6475102e-016 u0_mc=0.000636738                vsat_mc=1479.59                    lvsat_mc=-0.000577041 lu0_mc=-9.23262e-11               wvsat_mc=-0.000426122               pvsat_mc=1.66188e-10 wu0_mc=-1.14612e-10               pu0_mc=1.66188e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_18ud15_mac.30 nmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=0.39981866 k2=-0.048385059               cit=-0.00036223287             voff=-0.2349243 eta0=-0.70928395                etab=-0.0658                    u0=0.031 ua=-1.6723753e-009            ub=3.3460494e-018             uc=1.6668141e-010 vsat=83830.552                  a0=6.7696167                  ags=6.1222222 keta=0.02142678                 pclm=3.2803086                  pdiblc2=-0.058410575 agidl=1.1850999e-009             tvoff=-0.00247713                kt1=-0.27854464 kt2=-0.055802469               ute=-0.6                       ua1=3.8857372e-009 ub1=-2.2e-018                  uc1=-3.017284e-011             at=-15859.836 lvth0=6.5744939e-009             lk2=5.3554184e-009             lcit=3.5702377e-010 lvoff=2.2646047e-009             lua=3.4055723e-017             lub=-7.4827161e-026 luc=-1.3293805e-017            lvsat=0.0021260415               la0=-1.4814094e-006 lags=-3.3672222e-007            lketa=-2.0962331e-009            lpclm=-3.1614475e-007 lpdiblc2=1.1193473e-008             lagidl=-1.2279794e-016            ltvoff=3.88764e-010 lkt1=6.6538526e-009             lua1=-2.0228454e-016            luc1=7.3330617e-018 lat=0.0051295425               lu0=0                          lkt2=3.741358e-009 wvth0=-6.8216877e-009            wk2=4.9777715e-009             wcit=2.5063844e-010 wvoff=2.1401709e-008             weta0=2.5267556e-007             wetab=1.4688e-008 wua=4.9618818e-018             wub=-3.9342222e-025            wuc=-2.3200692e-017 wa0=-7.960496e-007             wags=-1.2355556e-006            wketa=-3.8228957e-008 wpclm=-7.7192889e-007            wpdiblc2=1.7197478e-008             wagidl=-1.5321349e-016 wtvoff=1.35408e-009               wkt1=1.9214203e-008             wua1=-4.5720499e-016 wub1=2.88e-025                  wuc1=3.712e-018                 pvth0=1.9821032e-016 pk2=-5.4673533e-016            pcit=-5.7222574e-017            pvoff=-8.638121e-016 pua=1.4124188e-023             pub=2.1550222e-032             puc=2.3201003e-024 pa0=1.8420591e-013             pags=5.3875556e-014             pketa=2.5693648e-015 ppclm=9.1049689e-014             ppdiblc2=-3.1403209e-015            pagidl=1.601081e-023 ptvoff=-1.16788e-016              pkt1=-1.6034163e-015            pua1=2.5205921e-023 puc1=-3.87904e-025              wat=0.0076227177               pat=-8.1427213e-010 wvsat=0.0070138425               pvsat=-1.0955939e-009            wu0=0 pu0=0                          leta0=6.6596173e-008             peta0=-1.9933956e-014 vsat_mc=-11530.9                   lvsat_mc=0.00130948                 wvsat_mc=0.00443555 pvsat_mc=-5.38755e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model pch_18ud15_mac.global pmos ( modelid=12                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=0                          igbmod=0 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_18ud15'          permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=3.65e-009                  toxm=3.65e-009                  dtox=4.74e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=1e-008 xw=0                          dlc=1.24e-008                  dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.43 k3=0.2                        k3b=0.4                        w0=0 dvt0=0.5                        dvt1=0.2                        dvt2=-0.09 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.4                       voffl=-5e-009 dvtp0=8e-007                     dvtp1=3                          lpe0=6e-008 lpeb=1e-007                     xj=8.5e-008                   ngate=1.15e+020 ndep=1e+017                     nsd=1e+020                     phin=0.15 cdsc=0                          cdscb=0                          cdscd=0 ud=0                          nfactor=0.8                        a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=1.2 delta=0.02                       pscbe1=9.264e+008                 pscbe2=1e-020 fprout=100                        pdits=0                          pditsd=0 pditsl=0                          rsh=16.7                       rdsw=200 prwg=0                          prwb=0                          wr=1 alpha0=0                          alpha1=0.055                      beta0=13.7 bgidl=9e+008                     cgidl=5                          egidl=0.5 aigbacc=0.01238                    bigbacc=0.006109                   cigbacc=0.2809 nigbacc=4.05                       aigbinv=0.35                       bigbinv=0.03 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1 aigc=0.009898                   bigc=0.001383                   cigc=1.515e-005 aigsd=0.0086                     bigsd=0.0004353                  cigsd=3.925e-020 nigc=1                          poxedge=1                          pigcd=1.672 ntox=1                          cgso=7.5e-012                   cgdo=7.5e-012 cgbo=0                          cgdl=1.105e-010                 cgsl=1.105e-010 clc=0                          cle=0.6                        cf='9.43e-011+5.68e-11*ccoflag_18ud15' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=5                          noff=2.6                        voffcv=-0.092 kt1l=0                          prt=0                          fnoimod=1 tnoimod=1                          em=7.46e+006                  ef=1.15 noia=0                          noib=0                          noic=0 lintnoi=-1.44e-008                 jss=2.81e-07                   jsd=2.81e-07 jsws=4.79e-14                   jswd=4.79e-14                   jswgs=4.79e-14 jswgd=4.79e-14                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=7.34                       bvd=7.34 xjbvs=1                          xjbvd=1                          jtssws=0 jtsswgs=5e-011                     jtsswgd=5e-011                     njtssw=20 njtsswg=8                          xtsswgs=0.46                       xtsswgd=0.46 tnjtsswg=1                          vtsswgs=7                          vtsswgd=7 pbs=0.830                      pbd=0.830                      cjs=0.001836 cjd=0.001836                   mjs=0.451                      mjd=0.451 pbsws=0.924                      pbswd=0.924                      cjsws=1.454e-010 cjswd=1.454e-010                 mjsws=0.560                      mjswd=0.560 pbswgs=0.949                      pbswgd=0.949                      cjswgs=1.847e-010 cjswgd=1.847e-010                 mjswgs=0.678                      mjswgd=0.678 tpb=0.00129                    tcj=0.00085                    tpbsw=0.00107 tcjsw=0.00066                    tpbswg=0.00140                    tcjswg=0.00100 xtis=3                          xtid=3                          dmcg=6.7e-008 dmci=6.7e-008                   dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=-5.1e-009 rshg=14.4                       gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          xrcrg1=12 xrcrg2=1                          pk2we=0                          lk2we=0 wk2we=0                          k2we=0                          pku0we=0 wku0we=-5e-10                     lku0we=0                          ku0we=0 pkvth0we=0                          wkvth0we=0                          lkvth0we=0 kvth0we=-0.005                     wec=-2800                      web=-150 scref=1e-6                       wpemod=1                          rnoia=0 rnoib=0                          tnoia=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.5 sigma_factor='sigma_factor_18ud15' ccoflag='ccoflag_18ud15' rcoflag='rcoflag_18ud15' rgflag='rgflag_18ud15' mismatchflag='mismatchflag_mos_18ud15' globalflag='globalflag_mos_18ud15' totalflag='totalflag_mos_18ud15' global_factor='global_factor_18ud15' local_factor='local_factor_18ud15' sigma_factor_flicker='sigma_factor_flicker_18ud15' noiseflag='noiseflagp_18ud15' noiseflag_mc='noiseflagp_18ud15_mc' delvto=0 mulu0=1 dlc_fmt=2 par1_io='par1_io' par2_io='par2_io' par3_io='par3_io' par4_io='par4_io' par5_io='par5_io' par6_io='par6_io' par7_io='par7_io' par8_io='par8_io' par9_io='par9_io' par10_io='par10_io' par11_io='par11_io' par12_io='par12_io' par13_io='par13_io' par14_io='par14_io' par15_io='par15_io' par16_io='par16_io' par17_io='par17_io' par18_io='par18_io' par19_io='par19_io' par20_io='par20_io' w7_io='2.0857*0.40825' w8_io='0.67082*0.40825' w9_io='0.54772*-0.10446' w10_io='0.54772*0.14211' w11_io='0.54772*-0.14894' w12_io='0.54772*0.78318' tox_c='toxp_18ud15'              dxl_c='dxlp_18ud15'              dxw_c='dxwp_18ud15' ddlc_c='ddlcp_18ud15'             cgo_c='cgop_18ud15'              cgl_c='cglp_18ud15' cj_c='cjp_18ud15'               cjsw_c='cjswp_18ud15'             cjswg_c='cjswgp_18ud15' cf_c='cfp_18ud15'               dvth_c='dvthp_18ud15'             dwvth_c='dwvthp_18ud15' dlvth_c='dlvthp_18ud15'            dpvth_c='dpvthp_18ud15'            du0_c='du0p_18ud15' dwu0_c='dwu0p_18ud15'             dlu0_c='dlu0p_18ud15'             dpu0_c='dpu0p_18ud15' dk2_c='dk2p_18ud15'              dwk2_c='dwk2p_18ud15'             dlk2_c='dlk2p_18ud15' dpk2_c='dpk2p_18ud15'             dags_c='dagsp_18ud15'             dwags_c='dwagsp_18ud15' dpdiblc2_c='dpdiblc2p_18ud15'         dlpdiblc2_c='dlpdiblc2p_18ud15'        dvsat_c='dvsatp_18ud15' dwvsat_c='dwvsatp_18ud15'           duc_c='ducp_18ud15'              dluc_c='dlucp_18ud15' dwuc_c='dwucp_18ud15'             dpuc_c='dpucp_18ud15'             dvoff_c='dvoffp_18ud15' dlvoff_c='dlvoffp_18ud15'           dwvoff_c='dwvoffp_18ud15'           dpvoff_c='dpvoffp_18ud15' dpkt1_c='dpkt1p_18ud15'            dltvoff_c='dltvoffp_18ud15'          dkt2_c='dkt2p_18ud15' duc1_c='duc1p_18ud15'             dlub1_c='dlub1p_18ud15'            dlketa_c='dlketap_18ud15' ss_flag_c='ss_flagp_18ud15'          ff_flag_c='ff_flagp_18ud15'          sf_flag_c='sf_flagp_18ud15' fs_flag_c='fs_flagp_18ud15'          monte_flag_c='monte_flagp_18ud15'      c1f_c='c1fp_18ud15' c2f_c='c2fp_18ud15'              c3f_c='c3fp_18ud15' global_mc='global_mc_flag_18ud15' tox_g='toxp_18ud15_ms_global'    dxl_g='dxlp_18ud15_ms_global' dxw_g='dxwp_18ud15_ms_global'    cgo_g='cgop_18ud15_ms_global' cgl_g='cglp_18ud15_ms_global'    cj_g='cjp_18ud15_ms_global' cjsw_g='cjswp_18ud15_ms_global'   cjswg_g='cjswgp_18ud15_ms_global' cf_g='cfp_18ud15_ms_global'     dvth_g='dvthp_18ud15_ms_global' dwvth_g='dwvthp_18ud15_ms_global'  dlvth_g='dlvthp_18ud15_ms_global' dpvth_g='dpvthp_18ud15_ms_global'  du0_g='du0p_18ud15_ms_global' dwu0_g='dwu0p_18ud15_ms_global'   dlu0_g='dlu0p_18ud15_ms_global' dpu0_g='dpu0p_18ud15_ms_global'   dk2_g='dk2p_18ud15_ms_global' dwk2_g='dwk2p_18ud15_ms_global'   dlk2_g='dlk2p_18ud15_ms_global' dpk2_g='dpk2p_18ud15_ms_global'   dags_g='dagsp_18ud15_ms_global' dwags_g='dwagsp_18ud15_ms_global'  dvsat_g='dvsatp_18ud15_ms_global' dwvsat_g='dwvsatp_18ud15_ms_global' dluc_g='dlucp_18ud15_ms_global' dlketa_g='dlketap_18ud15_ms_global' ss_flag_g='ss_flagp_18ud15_ms_global' ff_flag_g='ff_flagp_18ud15_ms_global'                                        monte_flag_g='monte_flagp_18ud15_ms_global' sf_flag_g='sf_flagp_18ud15_ms_global'                                        fs_flag_g='fs_flagp_18ud15_ms_global' weight1=-2.2915882 weight2=1.8541176 weight3=1.0677647 weight4=-0.58823529 weight5=-0.40837059 tox_1=8.0597748e-012 tox_2=-2.813774e-011 tox_3=-2.6572367e-012 tox_4=9.4219297e-011 tox_5=7.1465402e-013 dxl_1=4.8370644e-010 dxl_2=-1.6886243e-009 dxl_3=-1.5947618e-010 dxl_4=-5.6546372e-009 dxl_5=4.2889837e-011 dxl_max=-1.5e-008 dxw_1=-2.1173527e-009 dxw_2=-9.4864039e-010 dxw_3=2.3732503e-010 dxw_4=-3.7265088e-025 dxw_5=-1.1765292e-008 dxw_max=-1.2e-008 cgo_1=-6.0687e-014 cgo_2=3.5716e-014 cgo_3=9.6404e-015 cgo_4=-1.0732e-029 cgo_5=8.2291e-015 cgl_1=-8.9412e-013 cgl_2=5.2622e-013 cgl_3=1.4203e-013 cgl_4=6.9896e-029 cgl_5=1.2124e-013 cj_1=1.4856e-005 cj_2=-8.7433e-006 cj_3=-2.36e-006 cj_4=-1.0173e-021 cj_5=-2.0145e-006 cjsw_1=1.1765e-012 cjsw_2=-6.9242e-013 cjsw_3=-1.8689e-013 cjsw_4=-3.002e-028 cjsw_5=-1.5954e-013 cjswg_1=1.4945e-012 cjswg_2=-8.7957e-013 cjswg_3=-2.3741e-013 cjswg_4=-1.1184e-028 cjswg_5=-2.0266e-013 cf_1=-7.6304e-013 cf_2=4.4907e-013 cf_3=1.2121e-013 cf_4=1.2335e-028 cf_5=1.0347e-013 dvth_1=-0.0058524 dvth_2=-0.0029508 dvth_3=0.00049632 dvth_4=8.846e-019 dvth_5=0.0012874 dwvth_1=-8.4283e-010 dwvth_2=2.6991e-010 dwvth_3=8.6161e-012 dwvth_4=-1.2127e-025 dwvth_5=1.3345e-010 dlvth_1=5.5107e-012 dlvth_2=1.4314e-011 dlvth_3=1.5798e-013 dlvth_4=-5.104e-027 dlvth_5=-2.1038e-012 dpvth_1=-2.2752e-017 dpvth_2=-5.9246e-017 dpvth_3=1.037e-018 dpvth_4=3.3642e-032 dpvth_5=9.0017e-018 du0_1=4.9392e-005 du0_2=0.000151182 du0_3=5.45112e-006 du0_4=-1.18638e-020 du0_5=-2.10762e-005 dwu0_1=2.448595e-011 dwu0_2=4.523955e-011 dwu0_3=5.068635e-012 dwu0_4=-2.385185e-026 dwu0_5=-7.7231e-012 dlu0_1=-1.2014e-013 dlu0_2=5.4883e-014 dlu0_3=6.2137e-012 dlu0_4=4.8332e-028 dlu0_5=1.1889e-013 dpu0_1=1.4019e-018 dpu0_2=7.2864e-019 dpu0_3=-3.0081e-019 dpu0_4=-3.4041e-034 dpu0_5=-3.1086e-019 dk2_1=0.001956 dk2_2=0.0019536 dk2_3=4.0495e-005 dk2_4=5.3353e-019 dk2_5=-0.00049273 dwk2_1=1.1028e-010 dwk2_2=-6.4946e-011 dwk2_3=-5.1324e-013 dwk2_4=-1.4238e-026 dwk2_5=-1.4672e-011 dlk2_1=6.5058e-012 dlk2_2=-3.8103e-012 dlk2_3=-8.3213e-012 dlk2_4=-7.7694e-028 dlk2_5=-1.0029e-012 dpk2_1=4.5083e-017 dpk2_2=1.0373e-017 dpk2_3=-5.8341e-018 dpk2_4=-1.167e-032 dpk2_5=-9.1161e-018 dags_1=0.0013833 dags_2=0.00067001 dags_3=0.0010512 dags_4=4.564e-019 dags_5=-0.00026225 dwags_1=-2.2845e-010 dwags_2=-1.1932e-009 dwags_3=8.2049e-010 dwags_4=4.7756e-025 dwags_5=1.8205e-010 dvsat_1=-503.13 dvsat_2=-851.2 dvsat_3=376 dvsat_4=-7.7169e-013 dvsat_5=183.45 dwvsat_1=1.3657e-005 dwvsat_2=0.00031499 dwvsat_3=0.00023774 dwvsat_4=1.1389e-019 dwvsat_5=-1.8382e-005 dluc_1=1.8332e-019 dluc_2=-1.0882e-019 dluc_3=3.3527e-019 dluc_4=-4.584e-035 dluc_5=-1.8823e-020 dlketa_1=-6.1108e-011 dlketa_2=3.6274e-011 dlketa_3=-1.1176e-010 dlketa_4=-4.4625e-026 dlketa_5=6.2745e-012 ss_flag_1=0.054487 ss_flag_2=-0.031757 ss_flag_3=-0.13012 ss_flag_4=7.1537e-017 ss_flag_5=-0.0094 ff_flag_1=-0.061108 ff_flag_2=0.036274 ff_flag_3=-0.11176 ff_flag_4=-2.9739e-017 ff_flag_5=0.0062745 monte_flag_1=0.0604875 monte_flag_2=-0.211162 monte_flag_3=-0.0199425 monte_flag_4=-0.707113 monte_flag_5=0.00536337 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.9998 b_4=-0.0002176                 c_4=0.0002609                  d_4=-0.001733 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=-0.0025                    mis_a_2=-0.042                     mis_a_3=-0.006 mis_b_1=0.0022                     mis_b_2=-0.1236                    mis_b_3=0.0477 mis_c_1=0.9692                     mis_c_2=0                          mis_c_3=0 mis_d_1=0.0008                     mis_d_2=0                          mis_d_3=0 mis_e_1=0.0051                     mis_e_2=0.0482                     mis_e_3=-0.0277 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=0                          xl0=1e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=60                         co_rsd=16.7                       bidirectionflag=1 designflag=1 cf0=9.43e-011                  cco=5.68e-11 noimod=6                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718                      tnoiamax=1e1 tnoiac1=4162131.0367               tnoiac2=-17357183.454              rnoiamax=0.001 rnoiac1=-0.022218                  rnoiac2=0.74858 saref0=0.468e-6            sbref0=0.468e-6 samax=10e-6               sbmax=10e-6 samin=0.135e-6            sbmin=0.135e-6 rllodflag=0                   lreflod=1e-6                llodref=1 lod_clamp=-1e90 wlod0=0 ku00=-0e-9               lku00=0e-16               wku00=-0e-15 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=-0.6 kvth00=-0e-10              lkvth00=-0.0e-16            wkvth00=-0e-16 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0.0                 lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=-8e-9              lku000=1e-16             wku000=-2.5e-15     		pku000=0 llodku000=1                   wlodku000=1 kvth000=-0e-10             lkvth000=-0.5e-16	      wkvth000=-3.5e-16     		pkvth000=0 llodvth00=1                   wlodvth00=1                  steta000=0 stk200=0.5                 lodk200=1 lodeta000=1 wlod1=0                   llod1=0.4e-6 ku01=-2.35e-7            lku01=15e-14              wku01=1e-14 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=-1 kvth01=0.5e-8              lkvth01=-15e-22             wkvth01=3e-15 pkvth01=0e-29               llodvth1=2                   wlodvth1=1 steta01=1                  lodeta01=1 stk21=-0.0                lodk21=1 wlod2=0 ku02=0                   lku02=0                   wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0 kvth02=0                   lkvth02=0                   wkvth02=0 pkvth02=0                   llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0       		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0                   lku03=0                   wku03=0 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0 kvth03=0                   lkvth03=0                   wkvth03=0 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=0e-2                lku003=-0e-9               wku003=0e-9        		pku003=0 llodku003=1                   wlodku003=1 kvth003=0.000               lkvth003=0.0e-10             wkvth003=0e-9       		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=4.68e-7             sa_b1=1.35e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.98e-7             spamax=16e-7               spamin=1.98e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc='2.0e-6*0'          ldpckvth0='0.6+0.4'           pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc='6.3e-4*0'          ldpcku0='0.5*2'             pku0dpc=0.0e-14 keta0dpc=-0.04               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc='0'                 wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='-0.000'            wkvth0dpl=0                   wdplkvth0=1 lkvth0dpl='-0.5e-7*0'         ldplkvth0='0.8+0.2'           pkvth0dpl=0 ku0dpl='1*0'               wku0dpl=0                   wdplku0=1 lku0dpl='1.70e-3'           ldplku0='0.5'               pku0dpl=-2e-11 keta0dpl=0.05                wketa0dpl=0                   wdplketa0=1 kvsatdpl=0.04                wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=0.0e-6              wkvth0dpx=0                   wdpxkvth0=1 lkvth0dpx=0e-10               ldpxkvth0=1                   pkvth0dpx=0 ku0dpx=0                   wku0dpx=0                   wdpxku0=1 lku0dpx=0                   ldpxku0=1                   pku0dpx=0 keta0dpx=0                   wketa0dpx=0                   wdpxketa0=1 kvsatdpx=0                   wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0.000              wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-10            ldpskvth0=1.0                 pkvth0dps=0 ku0dps=-0.01               wku0dps=0                   wdpsku0=1 lku0dps=0.0e-14             ldpsku0=1                   pku0dps=0 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=0.00                wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa=0.0e-9              ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa=-0.0                wku0dpa=0e-9                wdpaku0=1 lku0dpa=-0e-8               ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                   wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.31e-7             spbmax='16e-7+1.6e-6+0.135e-6'    spbmin='1.98e-7+0.198e-6+0.135e-6' pse_mode=1 kvth0dp2=0.0                 wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=5e-7                ldp2kvth0=0.6                 pkvth0dp2=0 ku0dp2=0.00                wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=2.5e-4              ldp2ku0=0.5                 pku0dp2=0 keta0dp2=-0.00               wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=-0.2                wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.0                wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0e-8               ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=1.0                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=10e-6               enxmax=10e-6		 enxmin=0.18e-6 kvth0enx='-0.025'            wkvth0enx='1e-9'              wenxkvth0=1.0 lkvth0enx='1e-7*0'            lenxkvth0=1.0                 pkvth0enx=-0e-17 ku0enx='-1.20+0.1'         wku0enx='-1.0e-7'           wenxku0=1.0 lku0enx='1e-11'             lenxku0=1.5                 pku0enx='-1.0e-15*0' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx='-0.5*0'            wka0enx=0                   wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx='-1*0'              wenx=0                   ku0enx0='0' eny0=8e-8 enyref=8e-8		 enymax=2.0e-6              enymin=0.045e-6 kvth0eny='-0.005*0'          wkvth0eny='-1.1e-8'           wenykvth0=1 lkvth0eny='1.0e-8*0'          lenykvth0=1.0                 pkvth0eny=0 ku0eny='1.1'               wku0eny='5.0e-7*1.2'        wenyku0=1 ku0eny0='-0.15'             wku0eny0='-1.0e-6*1'         weny0ku0=1 lku0eny='7.8e-7'            lenyku0='1.0'               pku0eny=-0.0e-16 keta0eny='0'                 wketa0eny=-5e-9               wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny='0'                 weny=1e-6 kvth0eny1='(-2.0e-4*0)'      wkvth0eny1='-1.0e-10*0'       weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1='(-8.0e-18)*0' ku0eny1='(-1e-2)*0.3'      wku0eny1='(-1.0e-10)*0'     weny1ku0=1 lku0eny1='(-1.0e-5)*0'      leny1ku0=1.0                pku0eny1='(-5.5e-17)*0' keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1='(1.0e-8)*0'       weny1ka0=1 lka0eny1='(4.0e-9)*0'       leny1ka0=1.0                pka0eny1='(3.0e-15)*0' kvsateny1=-0.0               weny1=1e-6 rx_mode=0 rxref=20e-6           ringxmax=9.027e-6            ringxmin=0.477e-6 kvth0rx='(0.02)*1'          wkvth0rx=-0.0e-5             wrxkvth0=1.0 lkvth0rx='(1.0e-9)*0'        lrxkvth0=1.0                 pkvth0rx=0.0e-17 ku0rx='(1.00)*0.6'        wku0rx=0.0e-4              wrxku0=1.0 lku0rx='(1.0e-5)*0'        lrxku0=1.0                 pku0rx='-1.0e-14*0' keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx='-0.3'              wrx=0                   ku0rx0=0.5 ry_mode=0 ryref=1.008e-5            ringymax=9.027e-6            ringymin=0.477e-6 kvth0ry='0.01*0'            wkvth0ry='-0.0e-5+2e-5*0'    wrykvth0=1.0 lkvth0ry='(1.0e-8)*0'        lrykvth0='1.0+0'             pkvth0ry=0.0e-16 ku0ry='-0.1'              wku0ry='-4.0e-7'           wryku0=1.0 lku0ry='2.5e-5*1'          lryku0='0.8'               pku0ry='(-5.0e-16)*0' keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry='-3.0*0'            wry=1e-6 kvth0ry0='(-0.01)*0'         ku0ry0='-0.09' sfxref=1.89e-7           sfxmax=3e-6               minwodx=0.53e-6 sfxmin=1.89e-7 lrefodx=5e-8              lodxref=1                 wodx=1e-6 kvth0odxa=-0.50             lkvth0odxa=2.0e-13           lodxakvth0=2.0 wkvth0odxa=-1.0e-12          wodxakvth0=2.0               pkvth0odxa=0.0e-16 ku0odxa=4.00              lku0odxa=2.0e-20           lodxaku0=3.0 wku0odxa=-1.0e-12          wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.3 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=0.5               r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.065             lku0odx1a=1.0e-7            lodx1aku0=1.0 wku0odx1a=-1.0e-12          wodx1aku0=2.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-1.5e-4           lkvth0odx1b=0.0e-7            lodx1bkvth0=0.5 wkvth0odx1b=2.0e-16           wodx1bkvth0=2.0               pkvth0odx1b=0.0e-16 ku0odx1b=0.000             lku0odx1b=0.0e-6            lodx1bku0=0.5 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=8.1e-7 sfymin=2.61e-7           sfymax=1e-6              minwody=9e-7 wody=1e-6 kvth0odya=0                 lkvth0odya=0e-5              lodyakvth0=1.0 wkvth0odya=0e-7              wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=-0.5              lku0odya=3.0e-7            lodyaku0=1.0 wku0odya=2.5e-5            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=-0e-2             wketa0ody=0                 wodyketa0=1 kvsatody=-0.0 lrefody=5.0e-8            lodyref=0.5 kvth0odyb=-0.00             lkvth0odyb=3.0e-9            lodybkvth0=1.0 wkvth0odyb=1.0e-8            wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.00             lku0odyb=0.0e-10           lodybku0=1.0 wku0odyb=-0.0e-7           wodybku0=1.0               pku0odyb=-0e-16 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model pch_18ud15_mac.1 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-006                     wmax=0.00090001                 vth0=-0.401958 k2=0.012                      cit=0.001                      voff=-0.14036 eta0=0.01                       etab=-0.04                      u0=0.016 ua=1.79568e-009               ub=1.008e-018                 uc=3.9301875e-011 vsat=100000                     a0=1.9939049                  ags=0.6081735 keta=-0.04                      pclm=0.9                        pdiblc2=0.0009 agidl=4.7253673e-011             tvoff=0.0032832                  kt1=-0.168988 kt2=-0.041                     ute=-0.8                       ua1=3.1290656e-009 ub1=-3.6373047e-018            uc1=5.6e-011                   at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=0                          wk2=0                          wvoff=0 wu0=0                          wuc=0                          wags=0 pvth0=0                          pk2=0                          pvoff=0 pu0=0                          puc=0                          pkt1=0 wvsat=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18ud15_mac.2 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.40115041 k2=0.013223777                cit=0.00092040041              voff=-0.14001767 eta0=0.01                       etab=-0.04                      u0=0.015587121 ua=1.6651222e-009             ub=1.0503889e-018             uc=3.8167749e-011 vsat=100000                     a0=1.987791                   ags=0.57383228 keta=-0.038623737               pclm=0.81742424                 pdiblc2=0.00076237374 agidl=4.2750588e-011             tvoff=0.00322974                 kt1=-0.16566405 kt2=-0.041206439               ute=-0.8                       ua1=3.1444876e-009 ub1=-3.6425649e-018            uc1=5.820202e-011              at=120000 lvth0=-7.2763941e-009            lk2=-1.1026231e-008            lcit=7.171923e-010 lvoff=-3.0843826e-009            lu0=3.7200379e-009             lua=1.1763256e-015 lub=-3.8192389e-025            luc=1.0218479e-017             la0=5.5085825e-008 lags=3.0941442e-007             lketa=-1.2400126e-008            lpclm=7.4400758e-007 lpdiblc2=1.2400126e-009             lagidl=4.0572791e-017             ltvoff=4.81698e-010 lkt1=-2.9948785e-008            lkt2=1.8600189e-009             lua1=-1.3895213e-016 lub1=4.7393878e-026             luc1=-1.9840202e-017            wvth0=0 wk2=0                          wvoff=0                          wu0=0 wuc=0                          wags=0                          pvth0=0 pk2=0                          pvoff=0                          pu0=0 puc=0                          pkt1=0                          wvsat=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18ud15_mac.3 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.40892111 k2=0.011869991                cit=0.0021165083               voff=-0.13438143 eta0=0.01                       etab=-0.04                      u0=0.019 ua=3.2067129e-009             ub=3.4444444e-019             uc=1.5602944e-011 vsat=100000                     a0=1.9381799                  ags=0.56735612 keta=-0.045733333               pclm=1.5                        pdiblc2=0.0024688889 agidl=4.6131159e-011             tvoff=0.00478623                 kt1=-0.17221249 kt2=-0.036093778               ute=-1.0844444                 ua1=2.2689852e-009 ub1=-4.0072544e-018            uc1=-5.5111111e-012            at=134222.22 lvth0=1.1936711e-009             lk2=-9.5506042e-009            lcit=-5.8656533e-010 lvoff=-9.2278838e-009            lu0=0                          lua=-5.0400825e-016 lub=3.8755556e-025             luc=3.4814116e-017             la0=1.0916197e-007 lags=3.1647344e-007             lketa=-4.6506667e-009            lpdiblc2=-6.2008889e-010 lagidl=3.6887969e-017             ltvoff=-1.21488e-009              lkt1=-2.281099e-008 lkt2=-3.7127822e-009            lua1=8.1534545e-016             lub1=4.4490547e-025 luc1=4.9607111e-017             lute=3.1004444e-007             lat=-0.015502222 wvth0=0                          wk2=0                          wvoff=0 wu0=0                          wuc=0                          wags=0 pvth0=0                          pk2=0                          pvoff=0 pu0=0                          puc=0                          pkt1=0 wvsat=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18ud15_mac.4 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-006                     wmax=0.00090001                 vth0=-0.407056 k2=0.0095998443               cit=0.000732                   voff=-0.14001408 eta0=0.01                       etab=-0.04                      u0=0.019 ua=2.9915328e-009             ub=5.56256e-019               uc=2.437e-011 vsat=99809.68                   a0=2.5734947                  ags=0.55202753 keta=-0.0419357                 pclm=1.8588                     pdiblc2=0.00072 agidl=8.4252575e-011             tvoff=0.0034947                  kt1=-0.17739619 kt2=-0.0432912                 ute=-0.6                       ua1=3.779921e-009 ub1=-3.7095711e-018            uc1=5.952e-011                 at=184505.6 lvth0=0                          lk2=-8.0977104e-009            lcit=2.9952e-010 lvoff=-5.6229888e-009            lu0=0                          lua=-3.6629299e-016 lub=2.5199616e-025             luc=2.92032e-017               la0=-2.974395e-007 lags=3.2628373e-007             lketa=-7.081152e-009             lpclm=-2.29632e-007 lpdiblc2=4.992e-010                 lagidl=1.2490263e-017             ltvoff=-3.88303e-010 lkt1=-1.9493422e-008            lkt2=8.93568e-010               lua1=-1.5165344e-016 lub1=2.5438818e-025             luc1=7.9872e-018                lat=-0.047683584 lvsat=0.0001218048               wvth0=0                          wk2=0 wvoff=0                          wu0=0                          wuc=0 wags=0                          pvth0=0                          pk2=0 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18ud15_mac.5 pmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=9e-006                     wmax=0.00090001                 vth0=-0.41077747 k2=-0.00014433861             cit=0.0012040816               voff=-0.16088473 eta0=0.01                       etab=-0.04                      u0=0.018408163 ua=2.711669e-009              ub=7.4692245e-019             uc=4.1122449e-012 vsat=103343.29                  a0=2.7049935                  ags=1.0268346 keta=-0.063106429               pclm=1.6665306                  pdiblc2=0.0014081633 agidl=1.0241774e-010             tvoff=0.00249808                 kt1=-0.20564755 kt2=-0.047510204               ute=-0.6                       ua1=3.661101e-009 ub1=-3.3741003e-018            uc1=1.2261225e-010             at=100859.82 lvth0=1.4513731e-009             lk2=-4.297479e-009             lcit=1.1540816e-010 lvoff=2.5165627e-009             lu0=2.3081633e-010             lua=-2.5714611e-016 lub=1.7763624e-025             luc=3.7103725e-017             la0=-3.4872406e-007 lags=1.4110899e-007             lketa=1.1754321e-009             lpclm=-1.5464694e-007 lpdiblc2=2.3081633e-010             lagidl=5.4058472e-018             ltvoff=3.79455e-013 lkt1=-8.4753888e-009            lkt2=2.5389796e-009             lua1=-1.0531364e-016 lub1=1.2355454e-025             luc1=-1.6618775e-017            lat=-0.01506173 lvsat=-0.0012563031              wvth0=0                          wk2=0 wvoff=0                          wu0=0                          wuc=0 wags=0                          pvth0=0                          pk2=0 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          pvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18ud15_mac.6 pmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=9e-006                     wmax=0.00090001                 vth0=-0.39758914 k2=-0.0026614722              cit=-0.00074065983             voff=-0.15624747 eta0=-0.080308642               etab=-0.04                      u0=0.02 ua=1.2076376e-009             ub=1.1058111e-018             uc=1.4876543e-011 vsat=82498.122                  pvsat=0                          a0=0.81604938 ags=2                          keta=-0.067901235               pclm=0.78061728 pdiblc2=0.00041975309              agidl=2.1326999e-010             tvoff=0.00224107 kt1=-0.2156344                 kt2=-0.024839506               ute=-0.6 ua1=3.7437551e-009             ub1=-3.2771858e-018            uc1=-9.5209877e-011 at=-31701.184                 lvth0=-4.6093531e-010            lk2=-3.9324946e-009 lcit=3.9739568e-010             lvoff=1.8441603e-009             lu0=0 lua=-3.9061556e-017            lub=1.2559739e-025             luc=3.5542901e-017 la0=-7.482716e-008             lketa=1.870679e-009              lpclm=-2.6189506e-008 lpdiblc2=3.741358e-010              lagidl=-1.0667729e-017            ltvoff=3.76467e-011 lkt1=-7.0272955e-009            lkt2=-7.482716e-010             lua1=-1.172985e-016 lub1=1.0950195e-025             luc1=1.4965432e-017             lat=0.0041596155 lvsat=0.0017662462               leta0=1.3094753e-008             wvth0=0 wk2=0                          wvoff=0                          wu0=0 wuc=0                          wags=0                          pvth0=0 pk2=0                          pvoff=0                          pu0=0 puc=0                          pkt1=0                          wvsat=0 voff_mc=-0.0167716                 u0_ss=-0.000516049               u0_fs=-0.000516049 u0_sf=0.000516049                u0_mc=0.000645062                vsat_ss=5160.49 vsat_ff=5160.49                    vsat_mc=-7740.74                   pvsat_ss=0.0 pvsat_ff=0.0                        pvsat_mc=0.0                        lvoff_mc=2.43188e-09 lu0_ss=7.48272e-11                lu0_fs=7.48272e-11                lu0_sf=-7.48272e-11 lu0_mc=-9.3534e-11                lvsat_ss=-0.000748272               lvsat_ff=-0.000748272 lvsat_mc=0.00112241                 wvoff_mc=0.0                        wu0_ss=0.0 wu0_fs=0.0                        wu0_sf=0.0                        wu0_mc=0.0 pvoff_mc=0.0                        pu0_ss=0.0                        pu0_fs=0.0 pu0_sf=0.0                        pu0_mc=0.0                        wvsat_ss=0.0 wvsat_ff=0.0                        wvsat_mc=0.0 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_18ud15_mac.7 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-007                     wmax=9e-006                     vth0=-0.402012 k2=0.012074583                cit=0.001                      voff=-0.14063535 eta0=0.01                       etab=-0.04                      u0=0.016222222 ua=1.9158667e-009             ub=9.7666667e-019             uc=3.996e-011 vsat=100000                     a0=1.988877                   ags=0.60761164 keta=-0.040077569               pclm=0.92222222                 pdiblc2=0.00092103125 agidl=4.7240065e-011             tvoff=0.00329244                 kt1=-0.16798667 kt2=-0.041717188               ute=-0.77777778                ua1=3.2659211e-009 ub1=-3.7617004e-018            uc1=6.3111111e-011             at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=4.86e-010                  wk2=-6.7125e-010               wvoff=2.478123e-009 wu0=-2e-009                    wua=-1.08168e-015              wub=2.82e-025 wuc=-5.923125e-018             wa0=4.525035e-008              wags=5.056748e-009 wketa=6.98125e-010               wpclm=-2e-007                    wpdiblc2=-1.8928125e-010 wagidl=1.224697e-019              wtvoff=-8.32e-011                 wkt1=-9.012e-009 wkt2=6.4546875e-009             wute=-2e-007                    wua1=-1.2316996e-015 wub1=1.1195615e-024             wuc1=-6.4e-017                  pvth0=0 pk2=0                          pvoff=0                          pu0=0 puc=0                          pkt1=0                          wvsat=0 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.8 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=9e-007                     wmax=9e-006                     vth0=-0.40116998 k2=0.013304416                cit=0.00091723845              voff=-0.14030825 eta0=0.01                       etab=-0.04                      u0=0.015811668 ua=1.7837055e-009             ub=1.0220924e-018             uc=3.9027926e-011 vsat=100000                     a0=1.9867391                  ags=0.57366749 keta=-0.038635523               pclm=0.84311771                 pdiblc2=0.00079547452 agidl=4.2736969e-011             tvoff=0.00323612                 kt1=-0.16448258 kt2=-0.041953518               ute=-0.77471942                ua1=3.2933411e-009 ub1=-3.7718775e-018            uc1=6.5988098e-011             at=120000 lvth0=-7.5866452e-009            lk2=-1.1080796e-008            lcit=7.4568159e-010 lvoff=-2.9471485e-009            lu0=3.6990954e-009             lua=1.1907721e-015 lub=-4.0928573e-025            luc=8.3979855e-018             la0=1.9263133e-008 lags=3.0583684e-007             lketa=-1.2992835e-008            lpclm=7.127317e-007 lpdiblc2=1.1312661e-009             lagidl=4.0572898e-017             ltvoff=5.07454e-010 lkt1=-3.1571824e-008            lkt2=2.1293342e-009             lua1=-2.4705421e-016 lub1=9.1694912e-026             luc1=-2.5921654e-017            lute=-2.7555836e-008 wvth0=1.7609318e-010             wk2=-7.257543e-010             wvoff=2.6152048e-009 wu0=-2.0209192e-009            wua=-1.0672495e-015            wub=2.5466852e-025 wuc=-7.741598e-018             wa0=9.4674171e-009             wags=1.4831395e-009 wketa=1.0607402e-010             wpclm=-2.3124116e-007            wpdiblc2=-2.9790708e-010 wagidl=1.2257653e-019             wtvoff=-5.74734e-011              wkt1=-1.0633237e-008 wkt2=6.7237038e-009             wute=-2.2752525e-007            wua1=-1.3396817e-015 wub1=1.1638133e-024             wuc1=-7.0074702e-017            pvth0=2.7922604e-015 pk2=4.9108375e-016             wcit=2.845767e-011              pcit=-2.5640361e-016 pvoff=-1.2351071e-015            pu0=1.8848192e-016             pua=-1.3001859e-022 pub=2.4625659e-031             puc=1.6384442e-023             pa0=3.2240422e-013 pags=3.2198213e-014             pketa=5.3343793e-015             ppclm=2.8148287e-013 ppdiblc2=9.7871872e-016             pagidl=-9.624978e-028             ptvoff=-2.31797e-016 pkt1=1.4607349e-014             pkt2=-2.4238372e-015            pute=2.4800252e-013 pua1=9.7291869e-022             pub1=-3.9870931e-031            puc1=5.4733068e-023 wvsat=0                          pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.9 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=9e-007                     wmax=9e-006                     vth0=-0.4099936 k2=0.011710643                cit=0.0021721589               voff=-0.13477664 eta0=0.01                       etab=-0.04                      u0=0.019339338 ua=3.3965975e-009             ub=2.4354437e-019             uc=1.3353216e-011 vsat=100000                     a0=1.8414663                  ags=0.55955418 keta=-0.046783704               pclm=1.4927333                  pdiblc2=0.0025882201 agidl=4.6117898e-011             tvoff=0.00478525                 kt1=-0.17377529 kt2=-0.036745867               ute=-1.0844444                 ua1=2.3578601e-009 ub1=-4.1670581e-018            uc1=-6.8028746e-012            at=135802.47 lvth0=2.0311012e-009             lk2=-9.3435828e-009            lcit=-6.2218169e-010 lvoff=-8.9766048e-009            lu0=-1.4606538e-010            lua=-5.6728016e-016 lub=4.393316e-025              luc=3.6383419e-017             la0=1.7761048e-007 lags=3.2122034e-007             lketa=-4.1113185e-009            lpclm=4.6506667e-009 lpdiblc2=-8.2282663e-010            lagidl=3.6887685e-017             ltvoff=-1.18109e-009 lkt1=-2.1442774e-008            lkt2=-3.5470053e-009            lua1=7.7262003e-016 lub1=5.2244183e-025             luc1=5.3420506e-017             lute=3.1004444e-007 lat=-0.017224691               wvth0=9.65236e-009               wk2=1.4341326e-009 wvoff=3.5568594e-009             wu0=-3.0540444e-009            wua=-1.7089613e-015 wub=9.0810062e-025             wuc=2.0247555e-017             wa0=8.7042228e-007 wags=7.0217399e-008             wketa=9.4533333e-009             wpclm=6.54e-008 wpdiblc2=-1.0739813e-009            wagidl=1.1935323e-019             wtvoff=8.86423e-012 wkt1=1.4065197e-008             wkt2=5.8688e-009                wua1=-7.998745e-016 wub1=1.4382335e-024             wuc1=1.1625871e-017             pvth0=-7.5368704e-015 pk2=-1.863193e-015             wcit=-5.00855e-010              pcit=3.205472e-016 pvoff=-2.2615107e-015            pu0=1.3145884e-015             pua=5.6944721e-022 pub=-4.659844e-031             puc=-1.4123736e-023            pa0=-6.1603658e-013 pags=-4.2722131e-014            pketa=-4.8541333e-015            ppclm=-4.1856e-014 ppdiblc2=1.8246397e-015             pagidl=2.5508907e-027             ptvoff=-3.04105e-016 pkt1=-1.2313945e-014            pkt2=-1.491992e-015             pua1=3.8452884e-022 pub1=-6.9782725e-031            puc1=-3.4320558e-023            wat=-0.014222222 pat=1.5502222e-008             wvsat=0                          pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.10 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=9e-007                     wmax=9e-006                     vth0=-0.40656669 k2=0.0099014634               cit=0.000760288                voff=-0.13928838 eta0=0.01                       etab=-0.04                      u0=0.019457778 ua=3.1571022e-009             ub=5.2890667e-019             uc=2.6751244e-011 vsat=98679.2                    a0=2.5804915                  ags=0.52853343 keta=-0.041804796               pclm=1.8986667                  pdiblc2=0.00024920373 agidl=8.4238763e-011             tvoff=0.00363514                 kt1=-0.17590903 kt2=-0.04377744                ute=-0.6                       ua1=3.8757364e-009 ub1=-3.7881719e-018            uc1=7.1125687e-011             at=178152.89 lvth0=-1.6212064e-010            lk2=-8.1857079e-009            lcit=2.8141568e-010 lvoff=-6.0890901e-009            lu0=-2.2186667e-010            lua=-4.140032e-016 lub=2.5669973e-025             luc=2.7808681e-017             la0=-2.9536567e-007 lags=3.4107362e-007             lketa=-7.2978192e-009            lpclm=-2.5514667e-007 lpdiblc2=6.7414388e-010             lagidl=1.2490331e-017             ltvoff=-4.4502e-010 lkt1=-2.0077177e-008            lkt2=9.532016e-010              lua1=-1.9882078e-016 lub1=2.7995466e-025             luc1=3.5462267e-018             lat=-0.04432896 lvsat=0.000845312                wvth0=-4.4038214e-009            wk2=-2.7145717e-009 wvoff=-6.5313e-009               wu0=-4.12e-009                 wua=-1.4901248e-015 wub=2.46144e-025               wuc=-2.14312e-017              wa0=-6.2971622e-008 wags=2.1144694e-007             wketa=-1.1781328e-009            wpclm=-3.588e-007 wpdiblc2=4.2371664e-009             wagidl=1.2430308e-019             wtvoff=-1.26389e-009 wkt1=-1.3384397e-008            wkt2=4.37616e-009               wua1=-8.6233891e-016 wub1=7.0740701e-025             wuc1=-1.0445119e-016            pvth0=1.4590857e-015 pk2=7.9197782e-016             wcit=-2.54592e-010              pcit=1.6293888e-016 pvoff=4.1949114e-015             pu0=1.9968e-015                pua=4.2939187e-022 pub=-4.233216e-032             puc=1.2550668e-023             pa0=-1.8664479e-014 pags=-1.3310903e-013            pketa=1.950005e-015              ppclm=2.29632e-013 ppdiblc2=-1.5744949e-015            pagidl=-6.170112e-028             ptvoff=5.10455e-016 pkt1=5.2537955e-015             pkt2=-5.367024e-016             pua1=4.2450606e-022 pub1=-2.3009831e-031            puc1=3.996876e-023              wat=0.0571744 pat=-3.0191616e-008            wvsat=0.01017432                 pvsat=-6.5115648e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.11 pmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=9e-007                     wmax=9e-006                     vth0=-0.41097908 k2=-0.00021865302             cit=0.0011620644               voff=-0.16155424 eta0=0.01                       etab=-0.04                      u0=0.018560091 ua=2.8051365e-009             ub=7.3100227e-019             uc=3.5260771e-012 vsat=105162.39                  a0=2.7640517                  ags=1.0169229 keta=-0.062722547               pclm=1.6357143                  pdiblc2=0.001392517 agidl=1.0240237e-010             tvoff=0.00248896                 kt1=-0.20512477 kt2=-0.048176446               ute=-0.6                       ua1=3.6664154e-009 ub1=-3.4087997e-018            uc1=1.2887769e-010             at=103169.81 lvth0=1.5587135e-009             lk2=-4.2388625e-009            lcit=1.2472288e-010 lvoff=2.5945967e-009             lu0=1.2823129e-010             lua=-2.7673658e-016 lub=1.7788245e-025             luc=3.6866497e-017             la0=-3.6695417e-007 lags=1.5060174e-007             lketa=8.6010351e-010             lpclm=-1.5259524e-007 lpdiblc2=2.282517e-010              lagidl=5.4065252e-018             ltvoff=1.98752e-012 lkt1=-8.6830372e-009            lkt2=2.6688138e-009             lua1=-1.1718558e-016 lub1=1.319995e-025              luc1=-1.8977054e-017            lat=-0.01508556 lvsat=-0.0016831304              wvth0=1.8145117e-009             wk2=6.6882968e-010 wvoff=6.0256664e-009             wu0=-1.3673469e-009            wua=-8.4120777e-016 wub=1.4328163e-025             wuc=5.2755102e-018             wa0=-5.3152413e-007 wags=8.9205187e-008             wketa=-3.4549346e-009            wpclm=2.7734694e-007 wpdiblc2=1.4081633e-010             wagidl=1.3836739e-019             wtvoff=8.20817e-011 wkt1=-4.7050142e-009            wkt2=5.9961735e-009             wua1=-4.7829612e-017 wub1=3.1229507e-025             wuc1=-5.6389009e-017            pvth0=-9.6606419e-016 pk2=-5.2754874e-016            wcit=3.781551e-010              pcit=-8.383249e-017 pvoff=-7.0230553e-016            pu0=9.2326531e-016             pua=1.7631423e-022 pub=-2.2158367e-033            puc=2.135051e-024              pa0=1.64071e-013 pags=-8.5434752e-014            pketa=2.8379577e-015             ppclm=-1.8465306e-014 ppdiblc2=2.3081633e-017             pagidl=-6.1020912e-027            ptvoff=-1.44725e-017 pkt1=1.868836e-015              pkt2=-1.1685076e-015            pua1=1.0684743e-022 pub1=-7.6004654e-032            puc1=2.122451e-023              wat=-0.020789923 pat=2.1446984e-010             wvsat=-0.016371861               pvsat=3.841446e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.12 pmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=9e-007                     wmax=9e-006                     vth0=-0.39818946 k2=-0.001171445               cit=-0.00075657514             voff=-0.15795044 eta0=-0.081742113               etab=-0.04                      u0=0.019444444 ua=1.2923574e-009             ub=8.9500274e-019             uc=1.4087791e-011 vsat=77006.788                  a0=0.55005298                 ags=2.1989026 keta=-0.070012324               pclm=0.7840192                  pdiblc2=1.3717421e-005 agidl=2.1340005e-010             tvoff=0.00244298                 kt1=-0.21232993 kt2=-0.024879115               ute=-0.6                       ua1=3.6229919e-009 ub1=-3.3591543e-018            uc1=-1.1961965e-010            at=-26302.869 lvth0=-2.9578204e-010            lk2=-4.1007077e-009            lcit=4.0292562e-010 lvoff=2.0720454e-009             lu0=0                          lua=-5.7383599e-017 lub=1.5410238e-025             luc=3.5335048e-017             la0=-4.5924349e-008 lags=-2.0785322e-008            lketa=1.9171212e-009             lpclm=-2.9099451e-008 lpdiblc2=4.2817764e-010             lagidl=-1.0688139e-017            ltvoff=8.65508e-012 lkt1=-7.63829e-009              lkt2=-7.0929913e-010            lua1=-1.1088917e-016 lub1=1.2480092e-025             luc1=1.7055061e-017             lat=0.0036879787 lvsat=0.0023994312               leta0=1.3302606e-008             wvth0=5.4028927e-009 wk2=-1.3410245e-008            wvoff=1.5326774e-008             wu0=5e-009 wua=-7.6247784e-016            wub=1.8972753e-024             wuc=7.0987654e-018 wa0=2.3939676e-006             wags=-1.7901235e-006            wketa=1.8999807e-008 wpclm=-3.0617284e-008            wpdiblc2=3.654321e-009              wagidl=-1.1705527e-018 wtvoff=-1.81721e-009              wkt1=-2.9740288e-008            wkt2=3.5648148e-010 wua1=1.0868691e-015             wub1=7.3771646e-025             wuc1=2.19688e-016 pvth0=-1.4863794e-015            pk2=1.5139171e-015             wcit=1.4323781e-010 pcit=-4.9769483e-017            pvoff=-2.0509661e-015            pu0=0 pua=1.6489839e-022             pub=-2.5654492e-031            puc=1.870679e-024 pa0=-2.601253e-013             pags=1.870679e-013              pketa=-4.1797984e-016 ppclm=2.6189506e-014             ppdiblc2=-4.8637654e-016            pagidl=1.8369133e-025 ptvoff=2.60925e-016               pkt1=5.4989507e-015             pkt2=-3.5075231e-016 pua1=-5.7683884e-023            pub1=-1.3769076e-031            puc1=-1.8806656e-023 wat=-0.04858483                pat=4.2447314e-009             wvsat=0.049422007 pvsat=-5.6986649e-009            weta0=1.2901235e-008             peta0=-1.870679e-015 voff_mc=-0.0186351                 u0_ss=-0.000573388               u0_fs=-0.000573388 u0_sf=0.000573388                u0_mc=0.000716735                vsat_ss=4300.41 vsat_ff=5991.9                     vsat_mc=-8600.82                   lvoff_mc=2.70209e-09 lu0_ss=8.31413e-11                lu0_fs=8.31413e-11                lu0_sf=-8.31413e-11 lu0_mc=-1.03927e-10               lvsat_ss=-0.00062356                lvsat_ff=-0.000868827 lvsat_mc=0.00124712                 wvoff_mc=1.67716e-08                wu0_ss=5.16049e-10 wu0_fs=5.16049e-10                wu0_sf=-5.16049e-10               wu0_mc=-6.45062e-10 pvoff_mc=-2.43188e-15               pu0_ss=-7.48272e-17               pu0_fs=-7.48272e-17 pu0_sf=7.48272e-17                pu0_mc=9.3534e-17                 wvsat_ss=0.00774075 wvsat_ff=-0.00748271                wvsat_mc=0.00774074                 pvsat_ss=-1.12241e-09 pvsat_ff=1.08499e-09                pvsat_mc=-1.12241e-09 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.13 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.39531118 k2=0.011410214                cit=0.0009842875               voff=-0.13218809 eta0=-0.05                      etab=-0.04                      u0=0.011 ua=1.479e-010                 ub=1.5e-018                   uc=2.51775e-011 vsat=100000                     a0=1.9452161                  ags=0.59326045 keta=-0.034517813               pclm=1                          pdiblc2=0.00056239688 agidl=4.7282714e-011             tvoff=0.0032                     kt1=-0.184 kt2=-0.036863281               ute=-1                         ua1=8.6057278e-010 ub1=-1.016815e-018             uc1=5.9570313e-011             at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=-5.5447416e-009            wk2=-7.331769e-011             wvoff=-5.1244056e-009 wu0=2.7e-009                   wua=5.0949e-016                wub=-1.89e-025 wuc=7.381125e-018              wa0=8.4545167e-008             wags=1.7972821e-008 wketa=-4.3056562e-009            wpclm=-2.7e-007                  wpdiblc2=1.3348969e-010 wagidl=8.4085695e-020             wkt1=5.4e-009                   wkt2=2.0861719e-009 wua1=9.3311387e-016             wub1=-1.3508354e-024            wuc1=-6.0813281e-017 pvth0=0                          pk2=0                          wcit=1.414125e-011 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          weta0=5.4e-008 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.14 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.39419986 k2=0.012395738                cit=0.00091731156              voff=-0.13117562 eta0=-0.05                      etab=-0.04                      u0=0.010741263 ua=8.7658449e-011             ub=1.4715829e-018             uc=2.0112203e-011 vsat=100000                     a0=1.8757916                  ags=0.55103114 keta=-0.033841827               pclm=0.90125316                 pdiblc2=0.0002957318 agidl=4.2785948e-011             tvoff=0.00307951                 kt1=-0.18575143 kt2=-0.036909975               ute=-1.0275252                 ua1=7.5319206e-010 ub1=-8.7111413e-019            uc1=5.9802496e-011             at=120000 lvth0=-1.0012954e-008            lk2=-8.879572e-009             lcit=6.0345326e-010 lvoff=-9.1224027e-009            lu0=2.3312237e-009             lua=5.4277637e-016 lub=2.5603781e-025             luc=4.5638326e-017             la0=6.2551541e-007 lags=3.8048613e-007             lketa=-6.090632e-009             lpclm=8.8970906e-007 lpdiblc2=2.4026523e-009             lagidl=4.0515864e-017             ltvoff=1.08557e-009 lkt1=1.5780401e-008             lkt2=4.2071303e-010             lua1=9.6750026e-016 lub1=-1.3127651e-024            luc1=-2.0919764e-018            lute=2.4800252e-007 wvth0=-6.09701e-009              wk2=9.2056092e-011             wvoff=-5.6041638e-009 wu0=2.5424455e-009             wua=4.5919282e-016             wub=-1.4987296e-025 wuc=9.2825528e-018             wa0=1.0932018e-007             wags=2.1855857e-008 wketa=-4.208253e-009             wpclm=-2.8356307e-007            wpdiblc2=1.5186137e-010 wagidl=7.84955e-020               wtvoff=8.34744e-011               wkt1=8.5087296e-009 wkt2=2.1845157e-009             wua1=9.4645242e-016             wub1=-1.4468737e-024 wuc1=-6.4507661e-017            pvth0=4.9759387e-015             pk2=-1.4900178e-015 wcit=2.8391873e-011             pcit=-1.2839811e-016            pvoff=4.3226217e-015 pu0=1.4195665e-015             pua=4.5317756e-022             pub=-3.525346e-031 puc=-1.7131864e-023            pa0=-2.2322282e-013            pags=-3.4986149e-014 pketa=-8.7760344e-016            ppclm=1.2220324e-013             ppdiblc2=-1.655289e-016 pagidl=5.0367658e-026             ptvoff=-7.52104e-016              pkt1=-2.8009653e-014 pkt2=-8.8607815e-016            pua1=-1.2018033e-022            pub1=8.653047e-031 puc1=3.3286358e-023             wvsat=0                          weta0=5.4e-008 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.15 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.39996208 k2=0.014883551                cit=0.0020696064               voff=-0.1302703 eta0=-0.13533333                etab=-0.04                      u0=0.0098648889 ua=-1.9077493e-010            ub=2.2490293e-018             uc=4.1381726e-011 vsat=100000                     a0=3.2712492                  ags=0.69613197 keta=-0.028078298               pclm=1.6001667                  pdiblc2=0.0014439355 agidl=4.6047099e-011             tvoff=0.00713096                 kt1=-0.10423673 kt2=-0.028205644               ute=-1.0844444                 ua1=-9.6298657e-010 ub1=1.1255667e-019             uc1=1.402061e-010              at=120000 lvth0=-3.7321336e-009            lk2=-1.1591288e-008            lcit=-6.5254806e-010 lvoff=-1.0109198e-008            lu0=3.2864711e-009             lua=8.4626875e-016 lub=-5.9137877e-025            luc=2.2454545e-017             la0=-8.9553338e-007 lags=2.2232622e-007             lketa=-1.2372878e-008            lpclm=1.2789333e-007 lpdiblc2=1.1511103e-009             lagidl=3.6961209e-017             ltvoff=-3.33051e-009 lkt1=-7.3070624e-008            lkt2=-9.0670076e-009            lua1=2.838135e-015 lub1=-2.3849663e-024            luc1=-8.9731904e-017            lute=3.1004444e-007 leta0=9.3013333e-008             wvth0=6.2399706e-010             wk2=-1.4214846e-009 wvoff=-4.9884369e-010            wu0=5.47296e-009               wua=1.5196739e-015 wub=-8.9683584e-025            wuc=-4.9781039e-018            wa0=-4.1638232e-007 wags=-5.270261e-008             wketa=-7.3815313e-009            wpclm=-3.129e-008 wpdiblc2=-4.412519e-011             wagidl=1.8307159e-019             wtvoff=-2.10228e-009 wkt1=-4.8519503e-008            wkt2=-1.8174e-009               wua1=2.1888875e-015 wub1=-2.4134198e-024            wuc1=-1.206822e-016             pvth0=-2.3499591e-015 pk2=1.597416e-016              wcit=-4.0855771e-010            pcit=3.4787694e-016 pvoff=-1.2421772e-015            pu0=-1.7746944e-015            pua=-7.0274682e-022 pub=4.6165494e-031             puc=-1.5877486e-024            pa0=3.4979289e-013 pags=4.628258e-014              pketa=2.58127e-015               ppclm=-1.527744e-013 ppdiblc2=4.8096458e-017             pagidl=-6.3620283e-026            ptvoff=1.63037e-015 pkt1=3.415112e-014              pkt2=3.47601e-015               pua1=-1.4744346e-021 pub1=1.91884e-030               puc1=9.4516611e-023             wvsat=0 weta0=1.308e-007                 peta0=-8.3712e-014               pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.16 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.40768402 k2=0.0087845904               cit=9.528e-005                 voff=-0.14384124 eta0=0.01                       etab=-0.04                      u0=0.0072 ua=2.0966686e-010             ub=9.74e-019                  uc=-1.17636e-011 vsat=110920                     a0=1.6722643                  ags=0.68710533 keta=-0.031324387               pclm=3.438                      pdiblc2=0.004400916 agidl=8.4356068e-011             tvoff=0.00159134                 kt1=-0.19632062 kt2=-0.04617588                ute=-0.6                       ua1=2.5343215e-009 ub1=-4.2648589e-018            uc1=-1.5456797e-010            at=260554.48 lvth0=1.2099061e-009             lk2=-7.6879531e-009            lcit=6.110208e-010 lvoff=-1.4237958e-009            lu0=4.992e-009                 lua=5.8998601e-016 lub=2.2464e-025                luc=5.6467554e-017             la0=1.2781691e-007 lags=2.2810327e-007             lketa=-1.0295381e-008            lpclm=-1.04832e-006 lpdiblc2=-7.4135725e-010            lagidl=1.2443469e-017             ltvoff=2.14854e-010 lkt1=-1.4136933e-008            lkt2=2.4339432e-009             lua1=5.9985779e-016 lub1=4.1657968e-025             luc1=9.89235e-017               lat=-0.089954865 lvsat=-0.0069888                 wvth0=-3.3982229e-009            wk2=-1.709386e-009 wvoff=-2.4337246e-009            wu0=6.912e-009                 wua=1.162567e-015 wub=-1.5444e-025               wuc=1.323216e-017              wa0=7.5443284e-007 wags=6.8732222e-008             wketa=-1.0610501e-008            wpclm=-1.7442e-006 wpdiblc2=5.0062534e-010             wagidl=1.8728496e-020             wtvoff=5.75533e-010 wkt1=4.9860351e-009             wkt2=6.534756e-009              wua1=3.4493448e-016 wub1=1.1364253e-024             wuc1=9.8673103e-017             pvth0=2.2426171e-016 pk2=3.439985e-016              wcit=3.439152e-010              pcit=-1.3370573e-016 pvoff=-3.8534746e-018            pu0=-2.69568e-015              pua=-4.7419842e-022 pub=-1.34784e-032              puc=-1.3242317e-023            pa0=-3.9952881e-013 pags=-3.1435713e-014            pketa=4.6478106e-015             ppclm=9.43488e-013 ppdiblc2=-3.0054388e-016            pagidl=4.1559299e-026             ptvoff=-8.34321e-017 pkt1=-9.2424084e-017            pkt2=-1.8693698e-015            pua1=-2.9430465e-022 pub1=-3.5306084e-031            puc1=-4.5870786e-023            wat=-0.016987029 pat=1.0871699e-008             wvsat=-0.0008424                 pvsat=5.39136e-010 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.17 pmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.40753894 k2=0.0016329666               cit=0.0015803265               voff=-0.15398485 eta0=0.01                       etab=-0.04                      u0=0.017040816 ua=1.9633418e-009             ub=1.0368184e-018             uc=2.800949e-011 vsat=82890.709                  a0=2.2221681                  ags=1.0038749 keta=-0.072740356               pclm=0.75                       pdiblc2=0.0015826531 agidl=1.023909e-010              tvoff=0.00253363                 kt1=-0.20073526 kt2=-0.045133546               ute=-0.6                       ua1=3.9610468e-009 ub1=-3.4549351e-018            uc1=8.3762173e-011             at=63439.093 lvth0=1.1533251e-009             lk2=-4.8988198e-009            lcit=3.1852653e-011 lvoff=2.5322094e-009             lu0=1.1540816e-009             lua=-9.3947207e-017 lub=2.0014084e-025             luc=4.0956049e-017             la0=-8.6645564e-008 lags=1.0456314e-007             lketa=5.8568467e-009             lpclm=2.5871527e-022 lpdiblc2=3.5776531e-010             lagidl=5.4098825e-018             ltvoff=-1.52639e-010 lkt1=-1.2415225e-008            lkt2=2.0274329e-009             lua1=4.3434947e-017 lub1=1.0070942e-025             luc1=5.9747448e-018             lat=-0.013079865 lvsat=0.0039426237               wvth0=-1.2816169e-009            wk2=-9.9762799e-010 wvoff=-7.8679248e-010            wu0=0                          wua=-8.3592496e-017 wub=-1.3195286e-025            wuc=-1.6759561e-017            wa0=-4.3828852e-008 wags=1.0094838e-007             wketa=5.5610932e-009             wpclm=1.0744898e-006 wpdiblc2=-3.0306122e-011            wagidl=1.4868492e-019             wtvoff=4.18849e-011 wkt1=-8.6555782e-009            wkt2=3.2575638e-009             wua1=-3.1299786e-016 wub1=3.5381694e-025             wuc1=-1.5785043e-017            pvth0=-6.0121464e-016 pk2=6.6412865e-017             wcit=1.7191837e-012             pcit=-2.4928163e-019 pvoff=-6.46157e-016              pu0=0                          pua=1.1803797e-023 pub=-2.2248386e-032            puc=-1.5455461e-024            pa0=-8.8206748e-014 pags=-4.4000015e-014            pketa=-1.6591112e-015            ppclm=-1.5580102e-013 ppdiblc2=-9.3480612e-017            pagidl=-9.1237078e-027            ptvoff=1.24691e-016 pkt1=5.2278051e-015             pkt2=-5.9126487e-016            pua1=-3.7711039e-023 pub1=-4.7843583e-032            puc1=-1.2321092e-024            wat=0.014967725 pat=-1.5906554e-009            wvsat=0.003672648                pvsat=-1.2217327e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.18 pmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.38392 k2=-0.0039240909              cit=-0.00071423262             voff=-0.12808665 eta0=-0.10611111                etab=-0.04                      u0=0.025 ua=1.0287909e-010             ub=3.5578272e-018             uc=-4.6989506e-011 vsat=114786.71                  a0=3.2609657                  ags=0.82191358 keta=-0.044858145               pclm=0.94351852                 pdiblc2=0.01062963 agidl=2.1396888e-010             tvoff=-0.00504198                kt1=-0.38101063 kt2=-0.013479784               ute=-0.6                       ua1=6.3968329e-009 ub1=-1.2072543e-018            uc1=2.6734484e-010             at=-68335.812 lvth0=-2.2714205e-009            lk2=-4.0930465e-009            lcit=3.6456373e-010 lvoff=-1.2230284e-009            lu0=0                          lua=1.7581988e-016 lub=-1.6540544e-025            luc=5.1830903e-017             la0=-2.3727121e-007 lags=1.3094753e-007             lketa=1.8139261e-009             lpclm=-2.8060185e-008 lpdiblc2=-9.540463e-010             lagidl=-1.0768924e-017            ltvoff=9.45825e-010 lkt1=1.3724704e-008             lkt2=-2.5623626e-009            lua1=-3.0975405e-016 lub1=-2.252043e-025             luc1=-2.0644742e-017            lat=0.0060274959 lvsat=-0.00068229584             leta0=1.6836111e-008             wvth0=-7.4396159e-009 wk2=-1.0932864e-008            wvoff=-1.1550636e-008            wu0=0 wua=3.080526e-016              wub=-4.9926667e-025            wuc=6.2068333e-017 wa0=-4.58538e-008              wags=-5.5083333e-007            wketa=-3.6389544e-009 wpclm=-1.7416667e-007            wpdiblc2=-5.9e-009                  wagidl=-1.6824921e-018 wtvoff=4.91926e-009               wkt1=1.2207234e-007             wkt2=-9.9029167e-009 wua1=-1.4095878e-015            wub1=-1.1989936e-024            wuc1=-1.2858005e-016 pvth0=2.9169522e-016             pk2=1.5070221e-015             wcit=1.0512954e-010 pcit=-1.5243784e-017            pvoff=9.1460035e-016             pu0=0 pua=-4.4984742e-023            pub=3.1012117e-032             puc=-1.2975591e-023 pa0=-8.791313e-014             pags=5.0508333e-014             pketa=-3.2510426e-016 ppclm=2.5254167e-014             ppdiblc2=7.57625e-016               pagidl=2.5639697e-025 ptvoff=-5.82528e-016              pkt1=-1.3727744e-014            pkt2=1.3170048e-015 pua1=1.212945e-022              pub1=1.7731394e-031             puc1=1.5123167e-023 wat=-0.010755182               pat=2.139166e-009              wvsat=0.015420082 pvsat=-2.9251106e-009            weta0=3.4833333e-008             peta0=-5.0508333e-015 vsat_ss=5160.51                    vsat_ff=5805.55                    lvsat_ss=-0.000748274 lvsat_ff=-0.000841805               wvsat_ss=0.00696663                 wvsat_ff=-0.007315 pvsat_ss=-1.01016e-09               pvsat_ff=1.06068e-09 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.19 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.41310813 k2=0.013181082                cit=0.001031425                voff=-0.1515812 eta0=0.13                       etab=-0.035386                  u0=0.018 ua=1.8686e-009                ub=1.01e-018                  uc=6.053875e-011 vsat=100000                     a0=2.0978593                  ags=0.66021725 keta=-0.05947375                pclm=0.5                        pdiblc2=0.0004288 agidl=4.7195057e-011             tvoff=0.003                      kt1=-0.178 kt2=-0.02799                   ute=-1                         ua1=4.3441234e-009 ub1=-6.1777116e-018            uc1=-1.7997062e-010            at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=4.0656125e-009             wk2=-1.0295863e-009            wvoff=5.3478716e-009 wu0=-1.08e-009                 wua=-4.19688e-016              wub=7.56e-026 wuc=-1.171395e-017             wa0=2.1178692e-009             wags=-1.8183852e-008 wketa=9.17055e-009               wpdiblc2=2.05632e-010               wagidl=1.3142066e-019 wtvoff=1.08e-010                  wkt1=2.16e-009                  wkt2=-2.7054e-009 wua1=-9.4800347e-016            wub1=1.4360488e-024             wuc1=6.8538825e-017 pvth0=0                          pk2=0                          wcit=-1.1313e-011 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          weta0=-4.32e-008 wetab=-2.49156e-009              pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.20 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.41329725 k2=0.014715916                cit=0.00097129289              voff=-0.15207654 eta0=0.13                       etab=-0.035386                  u0=0.01689899 ua=1.5576555e-009             ub=1.1228535e-018             uc=5.9275782e-011 vsat=100000                     a0=1.9711439                  ags=0.6136996 keta=-0.059313123               pclm=0.40366162                 pdiblc2=0.00014374849 agidl=4.2679471e-011             tvoff=0.0030833                  kt1=-0.17124523 kt2=-0.028286997               ute=-1.0275252                 ua1=4.3396751e-009 ub1=-6.4988718e-018            uc1=-2.0025541e-010            at=120000 lvth0=1.7040278e-009             lk2=-1.3828852e-008            lcit=5.4179028e-010 lvoff=4.4630373e-009             lu0=9.920101e-009              lua=2.8016101e-015 lub=-1.0168103e-024            luc=1.1379344e-017             la0=1.1417053e-006 lags=4.1912405e-007             lketa=-1.4472497e-009            lpclm=8.6800884e-007 lpdiblc2=2.5683141e-009             lagidl=4.0685427e-017             ltvoff=-7.50518e-010 lkt1=-6.086044e-008             lkt2=2.6759473e-009             lua1=4.0078882e-017 lub1=2.8936534e-024             luc1=1.827659e-016              lute=2.4800252e-007 wvth0=4.2155827e-009             wk2=-1.1608397e-009            wvoff=5.6823351e-009 wu0=-7.8272727e-010            wua=-3.3460557e-016            wub=3.8440909e-026 wuc=-1.186578e-017             wa0=5.7829898e-008             wags=-1.1985114e-008 wketa=9.546247e-009              wpclm=-1.4863636e-008            wpdiblc2=2.3393236e-010 wagidl=1.3599296e-019             wtvoff=8.14313e-011               wkt1=6.7538284e-010 wkt2=-2.4718923e-009            wua1=-9.9024844e-016            wub1=1.5921155e-024 wuc1=7.5923608e-017             pvth0=-1.3512317e-015            pk2=1.1825935e-015 wcit=-7.5804941e-013            pcit=-9.5100105e-017            pvoff=-3.0135159e-015 pu0=-2.6784273e-015            pua=-7.6659267e-022            pub=3.3480341e-031 puc=1.3679858e-024             pa0=-5.0196538e-013            pags=-5.5850626e-014 pketa=-3.3850299e-015            ppclm=1.3392136e-013             ppdiblc2=-2.5498628e-016 pagidl=-4.1196354e-026            ptvoff=2.39384e-016               pkt1=1.3376401e-014 pkt2=-2.1039046e-015            pua1=3.8062721e-022             pub1=-1.4061613e-030 puc1=-6.6536894e-023            wvsat=0                          weta0=-4.32e-008 wetab=-2.49156e-009              pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.21 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.40721541 k2=0.015032352                cit=0.001980559                voff=-0.13947229 eta0=0.30066667                 etab=-0.035386                  u0=0.028844444 ua=5.6562395e-009             ub=-6.7755556e-019            uc=5.4562239e-011 vsat=100000                     a0=3.4160679                  ags=0.67369554 keta=-0.060365625               pclm=1.6266667                  pdiblc2=0.00091393778 agidl=4.629239e-011              tvoff=0.00221475                 kt1=-0.24681335 kt2=-0.024791644               ute=-1.6533333                 ua1=4.1195056e-009 ub1=-7.1906742e-018            uc1=-3.2069444e-010            at=120000 lvth0=-4.9251831e-009            lk2=-1.4173767e-008            lcit=-5.5830974e-010 lvoff=-9.2756027e-009            lu0=-3.1004444e-009            lua=-1.6658465e-015 lub=9.4563556e-025             luc=1.6517106e-017             la0=-4.3326184e-007 lags=3.5372847e-007             lketa=-3.0002226e-010            lpclm=-4.6506667e-007 lpdiblc2=1.7288078e-009             lagidl=3.6747345e-017             ltvoff=1.962e-010 lkt1=2.1508808e-008             lkt2=-1.1339876e-009            lua1=2.8006367e-016 lub1=3.647718e-024              luc1=3.1404444e-016             lute=9.3013333e-007 leta0=-1.8602667e-007            wvth0=4.5407943e-009             wk2=-1.501837e-009 wvoff=4.4702273e-009             wu0=-4.776e-009                wua=-1.6377139e-015 wub=6.8352e-025                wuc=-1.209558e-017             wa0=-4.9458445e-007 wags=-4.0586937e-008            wketa=1.0053625e-008             wpclm=-4.56e-008 wpdiblc2=2.420736e-010              wagidl=5.0614699e-020             wtvoff=5.52474e-010 wkt1=2.8471872e-008             wkt2=-3.66096e-009              wute=3.072e-007 wua1=-5.5565824e-016            wub1=1.5303248e-024             wuc1=1.2820409e-016 pvth0=-1.7057124e-015            pk2=1.5542806e-015             wcit=-3.6047213e-010 pcit=2.9698824e-016             pvoff=-1.6923184e-015            pu0=1.67424e-015 pua=6.5379541e-022             pub=-3.683328e-031             puc=1.6184687e-024 pa0=1.0016626e-013             pags=-2.4674639e-014            pketa=-3.938072e-015 ppclm=1.67424e-013               ppdiblc2=-2.6386022e-016            pagidl=5.1865946e-026 ptvoff=-2.74052e-016              pkt1=-1.6921773e-014            pkt2=-8.078208e-016 pute=-3.34848e-013              pua1=-9.3076108e-023            pub1=-1.3388095e-030 puc1=-1.2352262e-022            wvsat=0                          weta0=-1.0464e-007 peta0=6.69696e-014               wetab=-2.49156e-009              pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.22 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.41941866 k2=0.0039507069               cit=0.0002453415               voff=-0.15237506 eta0=0.01                       etab=-0.035386                  u0=0.024 ua=3.4130052e-009             ub=5.816e-019                 uc=7.3500742e-012 vsat=128080                     a0=4.6720865                  ags=1.1264257 keta=-0.06114159                pclm=-2.376                     pdiblc2=0.010191376 agidl=8.4051888e-011             tvoff=0.00199838                 kt1=-0.18593657 kt2=-0.02099976                ute=0.424                      ua1=6.2035499e-009 ub1=3.4545069e-019             uc1=3.104e-010                 at=188133.19 lvth0=2.8848948e-009             lk2=-7.0815148e-009            lcit=5.5222944e-010 lvoff=-1.0178299e-009            lu0=0                          lua=-2.3017653e-016 lub=1.39776e-025               luc=4.6732891e-017             la0=-1.2371137e-006 lags=6.3981186e-008             lketa=1.9659494e-010             lpclm=2.09664e-006 lpdiblc2=-4.2087528e-009            lagidl=1.2581267e-017             ltvoff=3.34678e-010 lkt1=-1.7452335e-008            lkt2=-3.5607936e-009            lua1=-1.0537247e-015 lub1=-1.1754019e-024            luc1=-8.9856e-017               lute=-3.9936e-007 lat=-0.043605242               lvsat=-0.0179712                 wvth0=2.9384815e-009 wk2=9.0091105e-010             wvoff=2.1745345e-009             wu0=-2.16e-009 wua=-5.6723569e-016            wub=5.7456e-026                wuc=2.9107759e-018 wa0=-8.6547115e-007            wags=-1.6850076e-007            wketa=5.4907883e-009 wpclm=1.39536e-006               wpdiblc2=-2.6262232e-009            wagidl=1.8298604e-019 wtvoff=3.55731e-010               wkt1=-6.2135649e-010            wkt2=-7.0603488e-009 wute=-5.5296e-007               wua1=-1.6364488e-015            wub1=-1.3531419e-024 wuc1=-1.524096e-016             pvth0=-6.802322e-016             pk2=1.6521823e-017 wcit=2.6288199e-010             pcit=-1.0195839e-016            pvoff=-2.2307507e-016 pu0=0                          pua=-3.1310647e-023            pub=3.234816e-032 puc=-7.9855994e-024            pa0=3.3753375e-013             pags=5.719021e-014 pketa=-1.0178564e-015            ppclm=-7.547904e-013             ppdiblc2=1.5718497e-015 pagidl=-3.2851713e-026            ptvoff=-1.48137e-016              pkt1=1.6978935e-015 pkt2=1.367788e-015              pute=2.156544e-013              pua1=5.9862987e-022 pub1=5.0660922e-031             puc1=5.6070144e-023             wat=0.022120465 pat=-1.4157098e-008            wvsat=-0.0101088                 pvsat=6.469632e-009 wetab=-2.49156e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.23 pmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.40677227 k2=-1.8126226e-005            cit=0.0018159699               voff=-0.16317012 eta0=0.01                       etab=-0.035386                  u0=0.017489796 ua=2.6017396e-009             ub=4.5126122e-019             uc=-1.2431551e-011 vsat=76245.946                  a0=2.7601536                  ags=1.0777029 keta=-0.054489395               pclm=4.6038776                  pdiblc2=-0.0035596574 agidl=1.0247858e-010             tvoff=0.00227369                 kt1=-0.2406208 kt2=-0.030018735               ute=-0.6                       ua1=3.7405818e-009 ub1=-2.5025679e-018            uc1=8.9469388e-011             at=99311.004 lvth0=-2.0471942e-009            lk2=-5.5336699e-009            lcit=-6.0315635e-011 lvoff=3.1922466e-009             lu0=2.5389796e-009             lua=8.6217053e-017 lub=1.9060812e-025             luc=5.4447725e-017             la0=-4.9145989e-007 lags=8.2983086e-008             lketa=-2.3977611e-009            lpclm=-6.2551225e-007 lpdiblc2=1.1541503e-009             lagidl=5.3948564e-018             ltvoff=2.27305e-010 lkt1=3.8745159e-009             lkt2=-4.3393469e-011            lua1=-9.3167113e-017 lub1=-6.4674649e-026            luc1=-3.6930612e-018            lat=-0.0089645894 lvsat=0.002244081                wvth0=-1.695616e-009             wk2=-1.0603785e-010 wvoff=4.1732576e-009             wu0=-2.4244898e-010            wua=-4.2832734e-016 wub=1.84248e-025               wuc=5.0786008e-018             wa0=-3.34341e-007 wags=6.1081273e-008             wketa=-4.2944258e-009            wpclm=-1.0066041e-006 wpdiblc2=2.7465415e-009             wagidl=1.0133957e-019             wtvoff=1.82248e-010 wkt1=1.2882614e-008             wkt2=-4.9044343e-009            wua1=-1.9394678e-016 wub1=-1.6046134e-025            wuc1=-1.8866939e-017            pvth0=1.1270658e-015 pk2=4.092319e-016              wcit=-1.2552823e-010            pcit=4.9521594e-017 pvoff=-1.0025771e-015            pu0=-7.478449e-016             pua=-8.5484904e-023 pub=-1.710072e-032             puc=-8.8310511e-024            pa0=1.3039299e-013 pags=-3.2346785e-014            pketa=2.798377e-015              ppclm=1.8197559e-013 ppdiblc2=-5.2352852e-016            pagidl=-1.0095906e-027            ptvoff=-8.04784e-017 pkt1=-3.568655e-015             pkt2=5.2698137e-016             pua1=3.6054074e-023 pub1=4.1463814e-032             puc1=3.9885061e-024             wat=-0.0044031077 pat=-3.8129044e-009            wvsat=0.0072608197               pvsat=-3.045197e-010 wetab=-2.49156e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.24 pmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=3.6e-007                   wmax=5.4e-007                   vth0=-0.47626 k2=-0.02690808                cit=-0.0017512325              voff=-0.17382284 eta0=-0.067407407               etab=-0.03538858                u0=0.055641975 ua=4.3955252e-009             ub=5.0318765e-018             uc=4.6904074e-010 vsat=157753.06                  a0=0.73309192                 ags=1.65 keta=-0.18204255                pclm=-1.6658272                 pdiblc2=0.0054320988 agidl=2.1318283e-010             tvoff=0.00970185                 kt1=0.087350273 kt2=-0.018237284               ute=-0.6                       ua1=2.2482457e-009 ub1=-3.5346902e-018            uc1=8.7741497e-011             at=52409.048 lvth0=8.0285259e-009             lk2=-1.6346267e-009            lcit=4.5692871e-010 lvoff=4.7368911e-009             lu0=-2.9930864e-009            lua=-1.7388186e-016 lub=-4.735811e-025             luc=-1.5365757e-017            la0=-1.9753595e-007 lags=6.9606132e-021             lketa=1.6097447e-008             lpclm=2.8359494e-007 lpdiblc2=-1.4965432e-010            lagidl=-1.065726e-017             ltvoff=-8.49778e-010 lkt1=-4.368129e-008             lkt2=-1.7517038e-009            lua1=1.2322163e-016 lub1=8.4983077e-026             luc1=-3.442517e-018             lat=-0.0021638056 lvsat=-0.0095744508              leta0=1.1224074e-008             wvth0=4.2423982e-008 wk2=1.4784898e-009             wvoff=1.3146907e-008             wu0=-1.6546667e-008 wua=-2.0099763e-015            wub=-1.2952533e-024            wuc=-2.16588e-016 wa0=1.319198e-006              wags=-9.98e-007                 wketa=7.0440625e-008 wpclm=1.23488e-006               wpdiblc2=-3.0933333e-009            wagidl=-1.2580287e-018 wtvoff=-3.04241e-009              wkt1=-1.3084254e-007            wkt2=-7.3338667e-009 wua1=8.3064933e-016             wub1=5.78218e-026               wuc1=-3.1594242e-017 pvth0=-5.2702759e-015            pk2=1.7947538e-016             wcit=6.6510948e-010 pcit=-6.5120875e-017            pvoff=-2.3037562e-015            pu0=1.6162667e-015 pua=1.438542e-022              pub=1.9742697e-031             puc=2.3310606e-023 pa0=-1.0937017e-013            pags=1.2122e-013                pketa=-8.0382053e-015 ppclm=-1.430396e-013             ppdiblc2=3.2325333e-016             pagidl=1.9609881e-025 ptvoff=3.87097e-016               pkt1=1.7271493e-014             pkt2=8.7924907e-016 pua1=-1.1251236e-022            pub1=9.812759e-033              puc1=5.833965e-024 wat=-0.075957406               pat=6.5624688e-009             wvsat=-0.0077817512 pvsat=1.8766531e-009             weta0=1.3933333e-008             peta0=-2.0203333e-015 wetab=-2.4901667e-009            letab=3.741358e-013              petab=-2.0203333e-019 u0_ss=-0.0020642                 vsat_ss=2580.26                    vsat_ff=-2580.22 vsat_fs=-25802.5                   lu0_ss=2.99309e-10                lvsat_ss=-0.000374134 lvsat_ff=0.000374134                lvsat_fs=0.00374136                 wu0_ss=1.11467e-09 pu0_ss=-1.61627e-16               wvsat_ss=0.00835997                 wvsat_ff=-0.00278667 wvsat_fs=0.0139333                  pvsat_ss=-1.2122e-09                pvsat_ff=4.04067e-10 pvsat_fs=-2.02033e-09 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.25 pmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.4072178 k2=0.010337252                cit=0.001                      voff=-0.1493905 eta0=0.01                       etab=-0.031111                  u0=0.011 ua=-1.868576e-010             ub=1.58e-018                  uc=1.5755e-011 vsat=100000                     a0=2.3196728                  ags=0.61152644 keta=-0.041525                  pclm=-1.1                       pdiblc2=0.00124 agidl=4.7193824e-011             tvoff=0.0026812                  kt1=-0.196 kt2=-0.041175                  ute=-1                         ua1=7.1821e-010 ub1=-1.0431195e-018            uc1=3.944625e-011              at=120000 lvth0=0                          lk2=0                          lvoff=0 lu0=0                          luc=0                          lketa=0 lpdiblc2=0                          ltvoff=0                          lub1=0 wvth0=1.9450944e-009             wk2=-5.80752e-012              wvoff=4.55922e-009 wu0=1.44e-009                  wua=3.2027674e-016             wub=-1.296e-025 wuc=4.4082e-018                wa0=-7.7735002e-008            wags=-6.5515968e-010 wketa=2.709e-009                 wpclm=5.76e-007                  wpdiblc2=-8.64e-011 wagidl=1.3186454e-019             wtvoff=2.22769e-010               wkt1=8.64e-009 wkt2=2.0412e-009                wua1=3.5732536e-016             wub1=-4.1240438e-025 wuc1=-1.045125e-017             pvth0=0                          pk2=0 pvoff=0                          pu0=0                          puc=0 pkt1=0                          wvsat=0                          wetab=-4.03056e-009 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.26 pmos ( level=54                         lmin=1.08e-006                  lmax=9e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.40853166 k2=0.011188961                cit=0.00097321277              voff=-0.15093456 eta0=0.01                       etab=-0.031111                  u0=0.010724748 ua=-3.0922078e-010            ub=1.6391793e-018             uc=1.6069992e-011 vsat=100000                     a0=2.2673298                  ags=0.56836068 keta=-0.042595044               pclm=-1.4578283                 pdiblc2=0.00094503939 agidl=4.2691464e-011             tvoff=0.00260815                 kt1=-0.19710407 kt2=-0.042413292               ute=-1.0275252                 ua1=5.4311156e-010 ub1=-7.9594151e-019            uc1=4.8032709e-011             at=120000 lvth0=1.1837875e-008             lk2=-7.6738936e-009            lcit=2.4135296e-010 lvoff=1.3911999e-008             lu0=2.4800252e-009             lua=1.1024922e-015 lub=-5.3320543e-025            luc=-2.8380789e-018            la0=4.7161053e-007 lags=3.8892346e-007             lketa=9.6410982e-009             lpclm=3.2240328e-006 lpdiblc2=2.6575951e-009             lagidl=4.0566257e-017             ltvoff=6.58202e-010 lkt1=9.9476913e-009             lkt2=1.1157014e-008             lua1=1.5776369e-015 lub1=-2.2270741e-024            luc1=-7.7364e-017               lute=2.4800252e-007 wvth0=2.4999686e-009             wk2=1.0886413e-010             wvoff=5.2712225e-009 wu0=1.44e-009                  wua=3.3746988e-016             wub=-1.4743636e-025 wuc=3.6883045e-018             wa0=-4.8797016e-008            wags=4.3368952e-009 wketa=3.5277386e-009             wpclm=6.5527273e-007             wpdiblc2=-5.4532364e-011 wagidl=1.3167534e-019             wtvoff=2.52486e-010               wkt1=9.9845646e-009 wkt2=2.6135739e-009             wua1=3.7651445e-016             wub1=-4.6093941e-025 wuc1=-1.3460115e-017            pvth0=-4.9994166e-015            pk2=-1.0331916e-015 wcit=-1.4492045e-012            pcit=1.3057333e-017             pvoff=-6.4151422e-015 pu0=-2.7655242e-029            pua=-1.5491023e-022            pub=1.6070564e-031 puc=6.486258e-024              pa0=-2.6073125e-013            pags=-4.4978415e-014 pketa=-7.3768351e-015            ppclm=-7.1424727e-013            ppdiblc2=-2.871274e-016 pagidl=1.7047297e-027             ptvoff=-2.67755e-016              pkt1=-1.2114527e-014 pkt2=-5.1570885e-015            pua1=-1.7289368e-022            pub1=4.3730063e-031 puc1=2.7109869e-023             wvsat=0                          wetab=-4.03056e-009 pvsat=0                          lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.27 pmos ( level=54                         lmin=6.3e-007                   lmax=1.08e-006 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.38154078 k2=0.011988572                cit=0.00093172194              voff=-0.12962813 eta0=0.01                       etab=-0.031111                  u0=0.0058888889 ua=-6.134567e-010             ub=1.3512729e-018             uc=-5.636298e-011 vsat=100000                     a0=3.98                       ags=1.1020547 keta=-0.030066444               pclm=1.5                        pdiblc2=0.0034844622 agidl=4.6059707e-011             tvoff=0.00312333                 kt1=-0.18733668 kt2=-0.038709056               ute=-0.8                       ua1=1.493459e-009 ub1=-3.1315556e-018            uc1=1.2949345e-010             at=120000 lvth0=-1.758218e-008             lk2=-8.5454701e-009            lcit=2.8657796e-010 lvoff=-9.3120175e-009            lu0=7.7511111e-009             lua=1.4341094e-015 lub=-2.1938745e-025            luc=7.6113861e-017             la0=-1.3952e-006 lags=-1.92803e-007              lketa=-4.0150756e-009            lpdiblc2=-1.1037582e-010 lagidl=3.6894873e-017             ltvoff=9.66513e-011               lkt1=-6.9876267e-010 lkt2=7.1193956e-009             lua1=5.4175819e-016             lub1=3.1874522e-025 luc1=-1.6615621e-016            wvth0=-4.702071e-009             wk2=-4.0607631e-010 wvoff=9.2632973e-010             wu0=3.488e-009                 wua=6.1937674e-016 wub=-4.685824e-026             wuc=2.7837498e-017             wa0=-6.976e-007 wags=-1.9479623e-007            wketa=-8.5408e-010               wpdiblc2=-6.833152e-010 wagidl=1.3438066e-019             wtvoff=2.25386e-010               wkt1=7.060272e-009 wkt2=1.349308e-009              wua1=3.8971854e-016             wub1=6.904214e-026 wuc1=-3.3863555e-017            pvth0=2.8508066e-015             pk2=-4.7190649e-016 wcit=1.71092e-011               pcit=-7.171328e-018             pvoff=-1.6792091e-015 pu0=-2.23232e-015              pua=-4.6218871e-022            pub=5.1075482e-032 puc=-1.9836363e-023            pa0=4.46464e-013               pags=1.7207669e-013 pketa=-2.6006528e-015            ppdiblc2=3.9824589e-016             pagidl=-1.2440719e-027 ptvoff=-2.38215e-016              pkt1=-8.9270477e-015            pkt2=-3.7790387e-015 pua1=-1.8728613e-022            pub1=-1.4037926e-031            puc1=4.9349619e-023 wvsat=0                          wetab=-4.03056e-009              pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.28 pmos ( level=54                         lmin=3.8e-007                   lmax=6.3e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.41019377 k2=0.0030112652               cit=0.0010100272               voff=-0.13574839 eta0=0.01                       etab=-0.031111                  u0=0.02424 ua=3.8688396e-009             ub=-1.794912e-019             uc=-4.4396586e-011 vsat=100000                     a0=2.6424                     ags=0.16970637 keta=-0.01205236                pclm=1.5                        pdiblc2=0.0039535594 agidl=8.4189551e-011             tvoff=0.00425066                 kt1=-0.20644631 kt2=-0.034075087               ute=-2.36                      ua1=-2.307265e-009 ub1=-3.8165232e-018            uc1=-5.702416e-010             at=247972.97 lvth0=7.557289e-010              lk2=-2.7999937e-009            lcit=2.3646256e-010 lvoff=-5.3950491e-009            lu0=-3.9936e-009               lua=-1.4345603e-015 lub=7.6030157e-025             luc=6.8455368e-017             la0=-5.39136e-007 lags=4.0389992e-007             lketa=-1.554409e-008             lpdiblc2=-4.1059799e-010 lagidl=1.2491773e-017             ltvoff=-6.24839e-010              lkt1=1.1531397e-008 lkt2=4.1536559e-009             lua1=2.9742215e-015             lub1=7.5712446e-025 luc1=2.8167422e-016             lute=9.984e-007                 lat=-0.081902698 wvth0=-3.8247875e-010            wk2=1.2391101e-009             wvoff=-3.8110656e-009 wu0=-2.2464e-009               wua=-7.3133609e-016            wub=3.3144883e-025 wuc=2.1539574e-017             wa0=-1.34784e-007              wags=1.7591819e-007 wketa=-1.2181334e-008            wpdiblc2=-3.806091e-010             wagidl=1.3342746e-019 wtvoff=-4.55089e-010              wkt1=6.7621511e-009             wkt2=-2.353231e-009 wute=4.4928e-007                wua1=1.4274445e-015             wub1=1.4516871e-025 wuc1=1.6462138e-016             pvth0=8.6267511e-017             pk2=-1.5248258e-015 wcit=-1.2404879e-011            pcit=1.1717683e-017             pvoff=1.3527238e-015 pu0=1.437696e-015              pua=4.022675e-022              pub=-1.9104104e-031 puc=-1.5805691e-023            pa0=8.626176e-014              pags=-6.5180536e-014 pketa=4.64879e-015               ppdiblc2=2.0451398e-016             pagidl=-6.3402394e-028 ptvoff=1.97289e-016               pkt1=-8.7362503e-015            pkt2=-1.4094138e-015 pute=-2.875392e-013             pua1=-8.5143076e-022            pub1=-1.8910027e-031 puc1=-7.7680737e-023            wat=0.00057814631              pat=-3.7001364e-010 wvsat=0                          wetab=-4.03056e-009              pvsat=0 lvsat=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.29 pmos ( level=54                         lmin=1.35e-007                  lmax=3.8e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.43056114 k2=0.0092244197               cit=0.0014678742               voff=-0.17816288 eta0=0.01                       etab=-0.031111                  u0=0.015183674 ua=1.0447253e-009             ub=9.8960408e-019             uc=9.0370204e-011 vsat=64593.959                  a0=-0.66702041                ags=1.4452466 keta=-0.082719775               pclm=1.855102                   pdiblc2=0.00059302106 agidl=1.0240033e-010             tvoff=0.000713536                kt1=-0.18769954 kt2=-0.015727666               ute=0.67346939                 ua1=6.4417772e-009 ub1=-1.6708538e-018            uc1=1.4050524e-010             at=192818.71 lvth0=8.6990057e-009             lk2=-5.223124e-009             lcit=5.7902235e-011 lvoff=1.1146601e-008             lu0=-4.6163265e-010            lua=-3.3315567e-016 lub=3.0435441e-025             luc=1.589632e-017              la0=7.5153796e-007 lags=-9.3560752e-008            lketa=1.2016202e-008             lpclm=-1.384898e-007 lpdiblc2=9.0001195e-010             lagidl=5.3895702e-018             ltvoff=7.54639e-010 lkt1=4.2201587e-009             lkt2=-3.0018384e-009            lua1=-4.3790491e-016 lub1=-7.9686595e-026            luc1=4.4829561e-018             lute=-1.8465306e-007 lat=-0.06039254                lvsat=0.013808356                wvth0=6.8683768e-009 wk2=-3.4333544e-009            wvoff=9.5706487e-009             wu0=5.877551e-010 wua=1.3219782e-016             wub=-9.5554286e-027            wuc=-3.1930031e-017 wa0=8.9944163e-007             wags=-7.1234461e-008            wketa=5.8685113e-009 wpclm=-1.7044898e-008            wpdiblc2=1.2515773e-009             wagidl=1.2951093e-019 wtvoff=7.43905e-010               wkt1=-6.1690383e-009            wkt2=-1.0049219e-008 wute=-4.5844898e-007            wua1=-1.1663771e-015            wub1=-4.5987843e-025 wuc1=-3.7239846e-017            pvth0=-2.7415662e-015            pk2=2.9743537e-016 wcit=-2.1379709e-013            pcit=6.9631606e-018             pvoff=-3.8661447e-015 pu0=3.3237551e-016             pua=6.5489276e-023             pub=-5.8049383e-032 puc=5.0474545e-024             pa0=-3.1708624e-013            pags=3.1208997e-014 pketa=-2.3906498e-015            ppclm=6.6475102e-015             ppdiblc2=-4.3203871e-016 pagidl=8.9342537e-028             ptvoff=-2.70319e-016              pkt1=-3.6930865e-015 pkt2=1.5920216e-015             pute=6.6475102e-014             pua1=1.6015968e-022 pub1=4.6868114e-032             puc1=1.0451399e-024             wat=-0.038065883 pat=1.4701158e-008             wvsat=0.011455535                pvsat=-4.4676587e-009 wetab=-4.03056e-009 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_18ud15_mac.30 pmos ( level=54                         lmin=9.45e-08                   lmax=1.35e-007 wmin=2.88e-07                   wmax=3.6e-007                   vth0=-0.17789498 k2=0.0045730355               cit=-0.0010313553              voff=-0.062123796 eta0=-0.18351852                etab=-0.03110713                u0=-0.039604938 ua=-9.1150672e-009            ub=-3.1629383e-019            uc=-1.0281975e-009 vsat=263689.69                  a0=12.847309                  ags=1.5740741 keta=0.18115642                 pclm=4.3059259                  pdiblc2=-0.016938272 agidl=2.1255226e-010             tvoff=0.00542245                 kt1=-0.085894107 kt2=-0.047860494               ute=-0.6                       ua1=7.6874158e-009 ub1=-6.8230429e-018            uc1=-1.2051585e-010            at=-760720.02 lvth0=-2.7937588e-008            lk2=-4.5486733e-009            lcit=4.2029051e-010 lvoff=-5.6790653e-009            lu0=7.482716e-009              lua=1.1400142e-015 lub=4.9370961e-025             luc=1.7808864e-016             la0=-1.2080398e-006 lags=-1.1224074e-007            lketa=-2.6245846e-008            lpclm=-4.9385926e-007 lpdiblc2=3.4420494e-009             lagidl=-1.058246e-017             ltvoff=7.1846e-011 lkt1=-1.0541629e-008            lkt2=1.6574216e-009             lua1=-6.1852251e-016 lub1=6.6738082e-025             luc1=4.2331014e-017             lat=0.077870577 lvsat=-0.015060524               leta0=2.8060185e-008             wvth0=-6.4987426e-008 wk2=-9.8547116e-009            wvoff=-2.706475e-008             wu0=1.7742222e-008 wua=2.8538369e-015             wub=6.30088e-025               wuc=3.2241778e-016 wa0=-3.0419201e-006            wags=-9.7066667e-007            wketa=-6.0311004e-008 wpclm=-9.1495111e-007            wpdiblc2=4.96e-009                  wagidl=-1.0310231e-018 wtvoff=-1.50183e-009              wkt1=-6.8474566e-008            wkt2=3.3304889e-009 wua1=-1.1274519e-015            wub1=1.2416288e-024             wuc1=4.3378402e-017 pvth0=7.6775253e-015             pk2=1.2285322e-015             wcit=4.0595367e-010 pcit=-5.1931122e-017            pvoff=1.4459881e-015             pu0=-2.1550222e-015 pua=-3.291484e-022             pub=-1.5079768e-031            puc=-4.6332978e-023 pa0=2.5441121e-013             pags=1.6162667e-013             pketa=7.2053799e-015 ppclm=1.3684391e-013             ppdiblc2=-9.6976e-016               pagidl=1.6917086e-025 ptvoff=5.53125e-017               pkt1=5.341215e-015              pkt2=-3.4803609e-016 pua1=1.5451552e-022             pub1=-1.9985043e-031            puc1=-1.0644506e-023 wat=0.21676906                 pat=-2.2249909e-008            wvsat=-0.045918936 pvsat=3.8516396e-009             weta0=5.5733333e-008             peta0=-8.0813333e-015 wetab=-4.0314889e-009            letab=-5.612037e-013             petab=1.3468889e-019 u0_ss=0.00516049                 vsat_ss=67086.1                    vsat_ff=-10320.9 vsat_fs=23222.2                    lu0_ss=-7.48272e-10               lvsat_ss=-0.00972754 lvsat_ff=0.00149655                 lvsat_fs=-0.00336723                wu0_ss=-1.48622e-09 pu0_ss=2.15502e-16                wvsat_ss=-0.0148623                 wvsat_ff=-2.2e-08 wvsat_fs=-0.00371558                pvsat_ss=2.15503e-09                pvsat_ff=2.2e-15 pvsat_fs=5.38758e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_hvt_mac.global nmos ( modelid=3                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_hvt'             permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=2.01e-009                  toxm=2.01e-009                  dtox=4.02e-010 epsrox=3.9                        wint=0                          lint=0 ll=0                          wl=0                          lln=1 wln=1                          lw=0                          ww=0 lwn=1                          wwn=1                          lwl=0 wwl=0                          llc=0                          wlc=0 lwc=0                          wwc=0                          lwlc=0 wwlc=0                          xl=-4e-009                    xw=6e-009 dlc=5.69006e-009               dwc=0                          xpart=1 toxref=3e-009                     dlcig=2.5e-009                   k1=0.48965 k3=-8.5                       k3b=2                          w0=0 dvt0=0.95                       dvt1=1.2                        dvt2=0.13 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.365                     voffl=0 dvtp0=1e-009                     dvtp1=0.7                        lpe0=1e-010 lpeb=1e-010                     xj=6.7e-008                   ngate=1.6e+020 ndep=1e+017                     nsd=1e+020                     phin=0.1404 cdsc=0                          cdscb=0                          cdscd=0 nfactor=1                          ud=0                          lud=0 wud=0                          pud=0                          a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=1                          drout=0.56                       pvag=2 delta=0.0075956                  pscbe1=1e+009                     pscbe2=1e-020 fprout=100                        pdits=0                          pditsd=0 pditsl=0                          rsh=18.0                       rdsw=120 rsw=100                        rdw=100                        prwg=0 prwb=0                          wr=1                          alpha0=2.772e-006 alpha1=1.8                        beta0=13.789                     agidl=1e-006 bgidl=2.388e+009                 cgidl=0.292                      egidl=0.27814 bigbacc=0.0021819                  cigbacc=0.25281                    nigbacc=4.05 aigbinv=0.2415                     bigbinv=0.0309                     cigbinv=0.006 eigbinv=1.1                        nigbinv=1                          cigc=0.00022705 cigsd=3.925e-020                 nigc=3.083                      poxedge=1 pigcd=3.5245                     ntox=1                          xrcrg1=12 xrcrg2=1                          vfbsdoff=0.01                       lvfbsdoff=0 wvfbsdoff=0                          pvfbsdoff=0                          cgso=6.81825e-011 cgdo=6.81825e-011               cgbo=0                          cgdl=2.91624e-011 cgsl=2.91624e-011               clc=0                          cle=0.6 cf='6.62e-11+9.73e-11*ccoflag_hvt'                                    ckappas=0.6 ckappad=0.6                        acde=0.4                        moin=5 noff=2.4373                     voffcv=-0.14                      tvfbsdoff=0.082 ltvfbsdoff=0                          wtvfbsdoff=0                          ptvfbsdoff=0 kt1l=0                          prt=0                          fnoimod=1 tnoimod=0                          em=1e+007                     ef=1.04 noia=0                          noib=0                          noic=0 lintnoi=-3.50e-008                 jss=2.2e-07                    jsd=2.2e-07 jsws=6.35e-14                   jswd=6.35e-14                   jswgs=6.35e-14 jswgd=6.35e-14                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=8.02                       bvd=8.02 xjbvs=1                          xjbvd=1                          njtsswg=4.12 xtsswgs=0.175                      xtsswgd=0.175                      tnjtsswg=1 vtsswgs=1                          vtsswgd=1                          pbs=0.748 pbd=0.748                      cjs=0.001686                   cjd=0.001686 mjs=0.406                      mjd=0.406                      pbsws=0.616 pbswd=0.616                      cjsws=1.31e-010                  cjswd=1.31e-010 mjsws=0.11                       mjswd=0.11                       pbswgs=0.944 pbswgd=0.944                      cjswgs=4.36e-010                  cjswgd=4.36e-010 mjswgs=0.7                        mjswgd=0.7                        tpb=0.00103 tcj=0.00075                    tpbsw=0.00067                    tcjsw=0.00016 tpbswg=0.0033                     tcjswg=0.00195                    xtis=3 xtid=3                          dmcg=3.8e-008                   dmci=3.8e-008 dmdg=0                          dmcgt=0                          dwj=0 xgw=0                          xgl=2.64e-009                  rshg=16.42 gbmin=1e-012                     rbpb=50                         rbpd=50 rbps=50                         rbdb=50                         rbsb=50 ngcon=1                          lnfactor=0                          pnfactor=0 wnfactor=0                          k2we=0                          ku0we=-0.0013 kvth0we=0.0005                     lk2we=0e-11                      lku0we=4.5e-11 lkvth0we=-1e-011                    pk2we=0e-18                      pku0we=-1e-18 pkvth0we=1.3e-018                   scref=1e-6                       web=2153.1 wec=-9093.6                    wk2we=0e-11                      wku0we=2e-11 wkvth0we=-4e-011                    wpemod=1 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.2                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.6 bidirectionflag='bidirectionflag_mos_hvt' iboffn_flag='iboffn_flag_hvt' iboffp_flag='iboffp_flag_hvt' sigma_factor='sigma_factor_hvt' ccoflag='ccoflag_hvt' rcoflag='rcoflag_hvt' rgflag='rgflag_hvt' mismatchflag='mismatchflag_mos_hvt' globalflag='globalflag_mos_hvt' totalflag='totalflag_mos_hvt' designflag='designflag_mos_hvt' global_factor='global_factor_hvt' local_factor='local_factor_hvt' sigma_factor_flicker='sigma_factor_flicker_hvt' noiseflag='noiseflagn_hvt' noiseflag_mc='noiseflagn_hvt_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w21='2.3875*0.35355' w22='0.70711*-0.35355' w23='0.54772*0.0088697' w24='0.54772*-0.21218' w25='0.54772*0.7283' w26='0.54772*-0.28609' w27='0.54772*-0.0042275' w28='0.54772*-0.30433' w29='0' w30='0' tox_c='toxn_hvt'                 ntox_c='ntoxn_hvt'                dxl_c='dxln_hvt' dxw_c='dxwn_hvt'                 cj_c='cjn_hvt'                  cjsw_c='cjswn_hvt' cjswg_c='cjswgn_hvt'               cgo_c='cgon_hvt'                 cgl_c='cgln_hvt' ddlc_c='ddlcn_hvt'                dvth_c='dvthn_hvt'                dlvth_c='dlvthn_hvt' dwvth_c='dwvthn_hvt'               dpvth_c='dpvthn_hvt'               du0_c='du0n_hvt' dlu0_c='dlu0n_hvt'                dwu0_c='dwu0n_hvt'                dpu0_c='dpu0n_hvt' dvsat_c='dvsatn_hvt'               dlvsat_c='dlvsatn_hvt'              dwvsat_c='dwvsatn_hvt' dpvsat_c='dpvsatn_hvt'              dvoff_c='dvoffn_hvt'               dlvoff_c='dlvoffn_hvt' dwvoff_c='dwvoffn_hvt'              dpvoff_c='dpvoffn_hvt'              dags_c='dagsn_hvt' dlags_c='dlagsn_hvt'               dwags_c='dwagsn_hvt'               dpags_c='dpagsn_hvt' dnfactor_c='dnfactorn_hvt'            dlnfactor_c='dlnfactorn_hvt'           dwnfactor_c='dwnfactorn_hvt' dpnfactor_c='dpnfactorn_hvt'           dcit_c='dcitn_hvt'                dlcit_c='dlcitn_hvt' dwcit_c='dwcitn_hvt'               dpcit_c='dpcitn_hvt'               deta0_c='deta0n_hvt' dleta0_c='dleta0n_hvt'              dweta0_c='dweta0n_hvt'              dpeta0_c='dpeta0n_hvt' dk2_c='dk2n_hvt'                 dlk2_c='dlk2n_hvt'                dpclm_c='dpclmn_hvt' dlpclm_c='dlpclmn_hvt'              dwpclm_c='dwpclmn_hvt'              dppclm_c='dppclmn_hvt' dua1_c='dua1n_hvt'                dlua1_c='dlua1n_hvt'               dwua1_c='dwua1n_hvt' dpua1_c='dpua1n_hvt'               dat_c='datn_hvt'                 dlat_c='dlatn_hvt' dwat_c='dwatn_hvt'                dpat_c='dpatn_hvt'                dkt1_c='dkt1n_hvt' dlkt1_c='dlkt1n_hvt'               dwkt1_c='dwkt1n_hvt'               dpkt1_c='dpkt1n_hvt' dkt2_c='dkt2n_hvt'                duc1_c='duc1n_hvt'                cf_c='cfn_hvt' jtsswg_c='jtsswgn_hvt'              dpdiblc2_c='dpdiblc2n_hvt'            dminv_c='dminvn_hvt' da0_c='da0n_hvt'                 ss_flag_c='ss_flagn_hvt'             ff_flag_c='ff_flagn_hvt' sf_flag_c='sf_flagn_hvt'             fs_flag_c='fs_flagn_hvt'             monte_flag_c='monte_flagn_hvt' c1f_c='c1fn_hvt'                 c2f_c='c2fn_hvt'                 c3f_c='c3fn_hvt' global_mc='global_mc_flag_hvt' tox_g='toxn_hvt_ms_global'       ntox_g='ntoxn_hvt_ms_global'      dxl_g='dxln_hvt_ms_global' dxw_g='dxwn_hvt_ms_global'       cj_g='cjn_hvt_ms_global'        cjsw_g='cjswn_hvt_ms_global' cjswg_g='cjswgn_hvt_ms_global'     cgo_g='cgon_hvt_ms_global'       cgl_g='cgln_hvt_ms_global' dvth_g='dvthn_hvt_ms_global'      dlvth_g='dlvthn_hvt_ms_global' dwvth_g='dwvthn_hvt_ms_global'     dpvth_g='dpvthn_hvt_ms_global'     du0_g='du0n_hvt_ms_global' dlu0_g='dlu0n_hvt_ms_global'      dwu0_g='dwu0n_hvt_ms_global'      dpu0_g='dpu0n_hvt_ms_global' dvsat_g='dvsatn_hvt_ms_global'     dlvsat_g='dlvsatn_hvt_ms_global' dwvsat_g='dwvsatn_hvt_ms_global'    dpvsat_g='dpvsatn_hvt_ms_global' dlvoff_g='dlvoffn_hvt_ms_global'    dags_g='dagsn_hvt_ms_global' dwags_g='dwagsn_hvt_ms_global'     deta0_g='deta0n_hvt_ms_global' dpeta0_g='dpeta0n_hvt_ms_global'    dk2_g='dk2n_hvt_ms_global'       dpclm_g='dpclmn_hvt_ms_global' dua1_g='dua1n_hvt_ms_global'      dlua1_g='dlua1n_hvt_ms_global' dpua1_g='dpua1n_hvt_ms_global'     dlat_g='dlatn_hvt_ms_global'      cf_g='cfn_hvt_ms_global' dpdiblc2_g='dpdiblc2n_hvt_ms_global'  dminv_g='dminvn_hvt_ms_global'     da0_g='da0n_hvt_ms_global' ss_flag_g='ss_flagn_hvt_ms_global'   ff_flag_g='ff_flagn_hvt_ms_global' monte_flag_g='monte_flagn_hvt_ms_global'                                       dpvoff_g='dpvoffn_hvt_ms_global' sf_flag_g='sf_flagn_hvt_ms_global'   fs_flag_g='fs_flagn_hvt_ms_global' weight1=-3.3752 weight2=1.9699333 weight3=-1.1658667 weight4=0.66666667 weight5=-0.46359333 tox_1=4.604223e-012 tox_2=-9.8935495e-012 tox_3=6.5248326e-013 tox_4=-3.7477187e-011 tox_5=8.6163431e-013 ntox_1=-0.0029406 ntox_2=0.00057423 ntox_3=-0.00037548 ntox_4=-1.3345e-018 ntox_5=0.00025595 dxl_1=1.0425052e-010 dxl_2=-2.2400112e-010 dxl_3=1.4773074e-011 dxl_4=8.4853424e-010 dxl_5=1.9509098e-011 dxl_max=-4e-009 dxw_1=-6.6805334e-010 dxw_2=-9.4440472e-010 dxw_3=-9.1243456e-011 dxw_4=3.2691163e-025 dxw_5=-5.8846294e-009 cj_1=1.1568e-005 cj_2=-2.259e-006 cj_3=1.4771e-006 cj_4=5.2498e-021 cj_5=-1.0069e-006 cjsw_1=8.9885e-013 cjsw_2=-1.7552e-013 cjsw_3=1.1477e-013 cjsw_4=-2.4513e-028 cjsw_5=-7.8235e-014 cjswg_1=2.9916e-012 cjswg_2=-5.8419e-013 cjswg_3=3.8199e-013 cjswg_4=1.9516e-027 cjswg_5=-2.6039e-013 cgo_1=-4.6783e-013 cgo_2=9.1356e-014 cgo_3=-5.9735e-014 cgo_4=9.2467e-028 cgo_5=4.072e-014 cgl_1=-2.001e-013 cgl_2=3.9074e-014 cgl_3=-2.555e-014 cgl_4=-2.5111e-028 cgl_5=1.7416e-014 dvth_1=0.0024119 dvth_2=0.0046204 dvth_3=-0.00099045 dvth_4=-2.0452e-018 dvth_5=-0.00090322 dlvth_1=1.1551e-010 dlvth_2=9.4689e-011 dlvth_3=6.494e-011 dlvth_4=2.5179e-025 dlvth_5=-2.6141e-011 dwvth_1=3.058e-010 dwvth_2=3.5355e-011 dwvth_3=-2.6486e-012 dwvth_4=4.128e-025 dwvth_5=-4.0851e-011 dpvth_1=1.6874e-017 dpvth_2=1.8183e-017 dpvth_3=6.2755e-019 dpvth_4=-2.2398e-032 dpvth_5=-4.1993e-018 du0_1=0.00032332 du0_2=0.00053619 du0_3=-5.9467e-005 du0_4=-1.4628e-019 du0_5=-0.00012925 dlu0_1=-2.7688e-012 dlu0_2=5.6312e-012 dlu0_3=3.9002e-012 dlu0_4=9.8483e-027 dlu0_5=-5.4583e-013 dwu0_1=-1.7645e-012 dwu0_2=3.768e-011 dwu0_3=-3.913e-012 dwu0_4=-3.0218e-027 dwu0_5=-5.0288e-012 dpu0_1=-1.8558e-019 dpu0_2=2.6352e-018 dpu0_3=-9.9627e-021 dpu0_4=1.3937e-033 dpu0_5=-5.3536e-019 dvsat_1=284.87 dvsat_2=4240.4 dvsat_3=-365.87 dvsat_4=-8.7648e-013 dvsat_5=-807.69 dlvsat_1=6.1692e-005 dlvsat_2=-1.2053e-005 dlvsat_3=4.4471e-005 dlvsat_4=-9.7672e-020 dlvsat_5=-5.9861e-006 dwvsat_1=3.7156e-005 dwvsat_2=0.0005523 dwvsat_3=-5.4984e-005 dwvsat_4=-6.7576e-020 dwvsat_5=-0.00010876 dwvsat_max=-0.002 dpvsat_1=8.845e-013 dpvsat_2=-1.7217e-013 dpvsat_3=-3.2941e-012 dpvsat_4=-8.6709e-028 dpvsat_5=-1.9591e-014 dlvoff_1=-9.5984e-012 dlvoff_2=1.8744e-012 dlvoff_3=-1.7303e-012 dlvoff_4=6.7338e-027 dlvoff_5=8.4394e-013 dags_1=0.076453 dags_2=0.069926 dags_3=-0.011037 dags_4=1.4282e-016 dags_5=-0.018223 dwags_1=1.4802e-010 dwags_2=-2.8843e-011 dwags_3=-3.7228e-010 dwags_4=-2.5184e-025 dwags_5=-6.294e-012 deta0_1=-6.8234e-005 deta0_2=1.3329e-005 deta0_3=-3.395e-005 deta0_4=-8.8272e-020 deta0_5=6.3642e-006 dpeta0_1=-9.8021e-019 dpeta0_2=1.9141e-019 dpeta0_3=-1.2516e-019 dpeta0_4=-2.3983e-033 dpeta0_5=8.5316e-020 dk2_1=0.00056814 dk2_2=0.001077 dk2_3=6.4015e-005 dk2_4=-1.5872e-018 dk2_5=-0.00021618 dpclm_1=-0.004901 dpclm_2=0.00095706 dpclm_3=-0.0006258 dpclm_4=-2.6081e-019 dpclm_5=0.00042658 dua1_1=1.7154e-011 dua1_2=-3.3497e-012 dua1_3=2.1903e-012 dua1_4=1.3138e-026 dua1_5=-1.493e-012 dlua1_1=-4.901e-019 dlua1_2=9.5706e-020 dlua1_3=-6.258e-020 dlua1_4=-3.7537e-034 dlua1_5=4.2658e-020 dpua1_1=-7.8416e-026 dpua1_2=1.5313e-026 dpua1_3=-1.0013e-026 dpua1_4=9.9218e-041 dpua1_5=6.8253e-027 dlat_1=3.2976e-005 dlat_2=-6.4538e-006 dlat_3=9.2541e-005 dlat_4=2.4741e-020 dlat_5=-4.3583e-006 cf_1=-4.5423e-013 cf_2=8.87e-014 cf_3=-5.7999e-014 cf_4=-8.9122e-028 cf_5=3.9536e-014 dpdiblc2_1=-4.901e-005 dpdiblc2_2=9.5706e-006 dpdiblc2_3=-6.258e-006 dpdiblc2_4=2.6992e-020 dpdiblc2_5=4.2658e-006 dminv_1=-0.0098021 dminv_2=0.0019141 dminv_3=-0.0012516 dminv_4=-7.0918e-018 dminv_5=0.00085316 da0_1=-0.017819 da0_2=0.0034725 da0_3=0.04189 da0_4=1.5018e-017 da0_5=0.00080694 ss_flag_1=0.047109 ss_flag_2=-0.0092197 ss_flag_3=0.1322 ss_flag_4=-1.659e-016 ss_flag_5=-0.0062261 ff_flag_1=-0.050911 ff_flag_2=0.0099215 ff_flag_3=0.11969 ff_flag_4=2.24e-017 ff_flag_5=0.0023055 monte_flag_1=0.086875 monte_flag_2=-0.186667 monte_flag_3=0.0123108 monte_flag_4=0.707108 monte_flag_5=0.0162575 sigma_local=1                          a_1=0.967413 b_1=-0.00234419                c_1=-0.00136694                d_1=0.000299617 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1.05039                    b_2=-0.00179548                c_2=-0.0041436 d_2=-0.000547178               a_3=1.01534                    b_3=-0.00514223 c_3=-0.0063604                 d_3=-0.00023778                e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.76 b_4=0.0009                     c_4=-0.007                     d_4=-1.0e-4 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=0.74                       b_5=-0.002                     c_5=-0.007 d_5=-1.0e-4                    e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.0025                     mis_a_2=0.047                      mis_a_3=0.1 mis_b_1=0.002                      mis_b_2=0                          mis_b_3=0 mis_c_1=0.1000                     mis_c_2=0.0000                     mis_c_3=0.0000 mis_d_1=0.00082                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.0063                     mis_e_2=0.0708                     mis_e_3=0.0368 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-4e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0 cf0=6.62e-11                   cco=9.73e-11 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.47                       l_rjtsswg=2.1e-5                     ll_rjtsswg=3 w_rjtsswg=0                          ww_rjtsswg=0                          p_rjtsswg=0.0 noimod=1                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6                sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=0                   lreflod=1e-6                llodref=3 lod_clamp=-1e90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=1 kvth00=0                   lkvth00=0                   wkvth00=0 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=0                   lku000=0                   wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0                   lkvth000=0                   wkvth000=0         		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=0                   wku01=0 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=0                   wkvth01=0 pkvth01=0                   llodvth1=1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.15               lku02=8e-7                wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=-0.5 kvth02=7e-3                lkvth02=-9e-9               wkvth02=16e-9 pkvth02=1e-15               llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=-0.03               lku03=7e5                 wku03=-5e-8 pku03=0                   tku03=0                   llodku03=-1 wlodku03=1                   kvsat3=0 kvth03=9e-3                lkvth03=-3e-9               wkvth03=-2e-8 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=-0.000                   lku003=-0.0e-9                   wku003=-0e-9         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0.0e-3                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='0.15*01'           wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl='1.4e-12*1'         ldplkvth0=1.5                 pkvth0dpl=0.0e-19 ku0dpl='0.50*0'            wku0dpl=0e-8                wdplku0=1 lku0dpl=5.0e-8              ldplku0=1.0                 pku0dpl=0.0e-11 keta0dpl='0.07*0'            wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0.00                wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx='0.25*1'            wku0dpx=0e-9                wdpxku0=1 lku0dpx='1.0e-8*1'          ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps='0.1*1'             wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='-0.70*1'           wku0dps=-0.0e-9             wdpsku0=1 lku0dps='9.0e-15*1'         ldpsku0=2.0                 pku0dps='-7.0e-23*0' keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps='-0.3*0'            wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa='0.01*0'            wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa='1.0e-9*0'          ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa='0.050*0'           wku0dpa=0e-7                wdpaku0=1 lku0dpa=0.0e-11             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=-0.0                wka0dpa=0                   wdpaka0=1 lka0dpa=-0.0e-7             ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa='1.5*0'             wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2='0.005*1'           wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2='3e-9*1'            ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.000               wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2='2.5e-5*1'          ldp2ku0=0.5                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2='0.5*0'             wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx='0.050*2'           wkvth0enx='8.0e-9*1'          wenxkvth0=1 lkvth0enx='1.0e-8*1'          lenxkvth0=1.0                 pkvth0enx=0 ku0enx='-0.90*1.0'         wku0enx='-0.9e-8*1.5'       wenxku0=1 lku0enx='2.0e-7*1'          lenxku0=1.0                 pku0enx='-3.0e-16*1.7' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0.0                 wka0enx=0                   wenxka0=1 lka0enx='1.0e-7*2'          lenxka0=1.0                 pka0enx='1.0e-14*1.7' kvsatenx=-0.0                wenx=0                   ku0enx0='0.15*0' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.01e-6 kvth0eny='0.04*1.7'          wkvth0eny='4.0e-10*4'         wenykvth0=1 lkvth0eny='1.0e-7*1.7'        lenykvth0=1.0                 pkvth0eny=0 ku0eny='-0.70*2'           wku0eny='-1.1e-8*1'         wenyku0=1 ku0eny0='0.025*0'           wku0eny0=0                   weny0ku0=1 lku0eny='6.0e-10*1.7'       lenyku0=1.5                 pku0eny=-0.0e-14 keta0eny=0.00                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-8             wenyka0=1 lka0eny='-6.0e-8*1.7'       lenyka0=1.0                 pka0eny='1.0e-14*1.7' kvsateny=-0.0                weny=0 kvth0eny1=0.000              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=0 ku0eny1='0.15*1.7'         wku0eny1=0.0e-8             weny1ku0=1 lku0eny1='1.0e-5*1.4'       leny1ku0=1.0                pku0eny1=-0.0e-14 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1.0                pka0eny1=0 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=-0.045              wkvth0rx=-0.0e-5             wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0.0e-16 ku0rx='0.3'               wku0rx=0.0e-8              wrxku0=1.0 lku0rx='-3.5e-10*0'        lrxku0=1                   pku0rx=0.0e-15 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.0                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=0.9027e-5           ringymin=0.117e-6 kvth0ry='-0.03*1'           wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry=0.0e-8              lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry='-0.02*1'           wku0ry=-0.0e-8             wryku0=1.0 lku0ry='-1.0e-8*1'         lryku0=1.0                 pku0ry=-0.0e-16 keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry=0                   wry=0 kvth0ry0=0.01                ku0ry0=0.02 sfxref=9.0e-8            sfxmax=3.906e-6           minwodx=0.0e-6 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0009            lkvth0odx1b=0.0e-7            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.0016           lku0odx1b=0.8e-10           lodx1bku0=1.0 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6              sfymax=10e-6             minwody=0.9e-6 wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-1.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.000            lkvth0odyb=0.0e-10           lodybkvth0=1.0 wkvth0odyb=-2.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.03             lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-1.0e-7           wodybku0=1.0               pku0odyb=0 web_mac=0  wec_mac=0 kvsatwe=0.0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_hvt_mac.1 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=9.01e-06                   vth0=0.62846448 lvth0=4.6445687e-012             wvth0=-2.6432436e-008            pvth0=-9.6231841e-019 k2=-0.051032045               lk2=1.9355542e-008             wk2=1.3152689e-009 pk2=-1.8275248e-014            cit=0.004                      voff=-0.20613951 lvoff=-4.4256733e-013            wvoff=-1.1171421e-008            pvoff=4.00966e-019 eta0=0.041125742                weta0=-1.6874923e-008            etab=-0.0072199256 wetab=-2.5187474e-009            u0=0.027441533                wu0=1.9945288e-009 ua=-1.3382438e-009            lua=3.3770637e-016             wua=2.3447228e-016 pua=-1.7264495e-022            ub=1.9096425e-018             lub=3.0608941e-031 wub=-3.8208016e-026            pub=-2.7566413e-036            uc=2.9401557e-010 luc=4.2574255e-017             wuc=2.3401576e-016             puc=-3.8342374e-022 vsat=130559.26                  wvsat=-0.0050366889              a0=0.46700304 la0=-8.9391377e-014            wa0=2.0056455e-008             pa0=-3.236798e-018 ags=2.2440312                  lags=1.7084405e-007             wags=-1.4205716e-006 pags=1.7997191e-012             keta=-0.24572293                lketa=-1.5834674e-008 wketa=2.6553214e-007             pketa=-1.6210053e-013            pclm=0.28881482 wpclm=1.0073378e-007             pdiblc2=0.00100058                 lpdiblc2=-5.2174332e-012 wpdiblc2=-5.2232329e-012            ppdiblc2=4.6988203e-017             aigbacc=0.010804139 laigbacc=-1.3797437e-009            waigbacc=-4.871472e-011             paigbacc=-9.9657995e-018 aigc=0.0098484605               laigc=-3.0375005e-012            waigc=1.9248664e-010 paigc=7.3535691e-017             bigc=0.0013527579               wbigc=1.3276712e-010 aigsd=0.0094385908               laigsd=7.4119488e-011             waigsd=4.8868809e-011 paigsd=-6.3657202e-017            bigsd=0.00057949723              wbigsd=4.5279833e-012 tvoff=0.00220302                 ltvoff=-2.89094e-010              wtvoff=-3.29911e-010 ptvoff=-2.81799e-018              kt1=-0.12875747                lkt1=-2.4664475e-012 wkt1=1.808193e-008              pkt1=-1.9486948e-018            kt2=-0.042975215 lkt2=-1.9144501e-015            wkt2=1.2078985e-008             pkt2=1.7241538e-020 ute=-0.678002                  wute=2.719812e-009              ua1=2.9095336e-009 lua1=-8.6390558e-023            wua1=-7.0754367e-016            pua1=-2.806762e-027 ub1=-2.0454315e-18             lub1=-2.2125973e-26             wub1=4.9715077e-25 pub1=2.0046134e-32              uc1=3.9624418e-010             luc1=-6.8349369e-016 wuc1=-4.0931474e-016            puc1=4.1987155e-022             at=153328.6 wat=-0.029977365               lcit=0                          wcit=0 pcit=0                          lu0=0                          pu0=0 lvsat=0                          pvsat=0                          lpclm=0 ppclm=0                          lat=0                          pat=0 leta0=0                          peta0=0                          jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=-0.000800517 voff_mc=-6.17113e-05               lvoff_mcl=5.19727e-09                lvoff_mc=5.55772e-10 wvoff_mcl=2.23698e-09                wvoff_mc=5.56389e-10                pvoff_mcl=-2.00434e-15 pvoff_mc=-5.01084e-15 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.2 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.61356386 lvth0=1.3355598e-008             wvth0=-1.4618826e-008            pvth0=-1.0585957e-014 k2=-0.02537011                lk2=-3.6375516e-009            wk2=-1.7114572e-008 pk2=-1.7621108e-015            cit=0.0048295845               voff=-0.19443738 lvoff=-1.0485555e-008            wvoff=-2.2291849e-008            pvoff=9.9643047e-015 eta0=0.041125742                weta0=-1.6874923e-008            etab=-0.0072199256 wetab=-2.5187474e-009            u0=0.027506294                wu0=4.0801523e-009 ua=-8.5328851e-010            lua=-9.6813563e-017            wua=2.6045515e-017 pua=1.4105431e-023             ub=1.9887574e-018             lub=-7.0886672e-026 wub=-5.9360938e-027            pub=-2.8918399e-032            uc=3.3686741e-010 luc=4.1790117e-018             wuc=-1.5190786e-016            puc=-3.7636179e-023 vsat=141024.66                  wvsat=-0.010028607               a0=0.90568107 la0=-3.9305561e-007            wa0=-3.7171783e-007            pa0=3.5102652e-013 ags=3.5273886                  lags=-9.7904423e-007            wags=-3.2671555e-007 pags=8.1962411e-013             keta=-0.23471794                lketa=-2.5695144e-008 wketa=2.2716586e-008             pketa=5.5462209e-014             pclm=0.26321898 wpclm=8.9128167e-008             pdiblc2=0.0010186384               lpdiblc2=-2.1397825e-011 wpdiblc2=-1.6785784e-010            ppdiblc2=1.9270881e-016             aigbacc=0.009648791 laigbacc=-3.445521e-010             waigbacc=-1.4974914e-011            paigbacc=-4.0196666e-017 aigc=0.010230824                laigc=-3.4563519e-010            waigc=2.8846584e-010 paigc=-1.246167e-017             bigc=0.0018499366               wbigc=6.7003587e-011 aigsd=0.0095390556               laigsd=-1.5897018e-011            waigsd=-5.7392714e-011 paigsd=3.1553122e-017             bigsd=0.00058012895              wbigsd=-1.161306e-012 tvoff=0.00197027                 ltvoff=-8.05463e-011              wtvoff=-6.30634e-010 ptvoff=2.6663e-016                kt1=-0.13734084                lkt1=7.6882394e-009 wkt1=1.810129e-008              pkt1=-1.9295482e-017            kt2=-0.049903879 lkt2=6.2080807e-009             wkt2=3.9389066e-008             pkt2=-2.4469815e-014 ute=-0.63873912                wute=-1.0403692e-008            ua1=2.84717e-009 lua1=5.5877691e-017             wua1=-2.7225063e-016            pua1=-3.9002537e-022 ub1=-1.3821062e-18             lub1=-6.1646545e-25             wub1=-1.9209013e-25 pub1=6.3760598e-31              uc1=-2.3818492e-010            luc1=-1.1504521e-016 wuc1=-3.9928069e-016            puc1=4.1088104e-022             at=151299.81 wat=-0.011706121               lcit=-7.4330767e-010            wcit=-3.3246176e-011 pcit=2.9788574e-017             lu0=-5.8025559e-011            pu0=-1.8687186e-015 lvsat=-0.0093769977              pvsat=4.4727588e-009             lpclm=2.2933864e-008 ppclm=1.0398627e-014             lbigc=-4.454721e-010             pbigc=5.8924125e-017 lbigsd=-5.6602301e-013            pbigsd=5.0976032e-018             lute=-3.5179541e-008 pute=1.1758659e-014             lat=0.001817792                pat=-1.6371034e-008 leta0=0                          peta0=0                          jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499997 voff_mc=0.00111217                 lvoff_mcl=-2.72e-15                  lvoff_mc=-4.9603e-10 wvoff_mcl=-3.91e-14                  wvoff_mc=-1.00274e-08               pvoff_mcl=-6e-21 pvoff_mc=4.4722e-15                 u0_ff=0.000220391                u0_ss=-0.000220391 u0_fs=0.000220391                u0_sf=-0.000220391               wu0_ff=-1.99674e-10 wu0_ss=1.99674e-10                wu0_fs=-1.99674e-10               wu0_sf=1.99674e-10 lu0_ff=-1.9747e-10                lu0_ss=1.9747e-10                 lu0_fs=-1.9747e-10 lu0_sf=1.9747e-10                 pu0_ff=1.78908e-16                pu0_ss=-1.78908e-16 pu0_fs=1.78908e-16                pu0_sf=-1.78908e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.3 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.66691341 lvth0=-1.0438301e-008            wvth0=-5.6511457e-008            pvth0=8.0981562e-015 k2=-0.022833783               lk2=-4.7687537e-009            wk2=-2.1411535e-008 pk2=1.5433455e-016             cit=0.0019919085               voff=-0.2304109 lvoff=5.558637e-009              wvoff=2.1496758e-008             pvoff=-9.5654137e-015 eta0=0.040897736                weta0=-1.4821503e-008            etab=-0.0072199256 wetab=-2.5187474e-009            u0=0.031761603                wu0=-1.4112113e-009 ua=-9.1531085e-010            lua=-6.9151597e-017            wua=3.2901325e-017 pua=1.104774e-023              ub=2.0745539e-018             lub=-1.0915188e-025 wub=-4.1991177e-026            pub=-1.2837832e-032            uc=5.7346362e-010 luc=-1.013429e-016             wuc=-3.2447382e-016            puc=3.932824e-023 vsat=115964.69                  wvsat=0.011864201                a0=0.094788613 la0=-3.139757e-008             wa0=1.1725487e-006             pa0=-3.3771633e-013 ags=1.3322222                  lags=0                          wags=1.5110067e-006 pags=0                          keta=-0.31953402                lketa=1.2132826e-008 wketa=1.7992603e-007             pketa=-1.46532e-014              pclm=0.11188431 wpclm=8.1700959e-008             pdiblc2=0.00094408086              lpdiblc2=1.1854857e-011 wpdiblc2=5.0360776e-010             ppdiblc2=-1.0676485e-016            aigbacc=0.0093885112 laigbacc=-2.2846728e-010            waigbacc=-1.6576067e-010            paigbacc=2.705378e-017 aigc=0.0090968476               laigc=1.6011827e-010             waigc=5.9151118e-010 paigc=-1.4761989e-016            bigc=0.00045109398              wbigc=5.7500571e-010 aigsd=0.0094900445               laigsd=5.9619427e-012             waigsd=1.8820481e-011 paigsd=-2.4379628e-018            bigsd=0.00057782687              wbigsd=1.95712e-011 tvoff=0.00217118                 ltvoff=-1.70151e-010              wtvoff=4.08252e-011 ptvoff=-3.28409e-017              kt1=-0.098165521               lkt1=-9.7839544e-009 wkt1=-5.0557817e-009            pkt1=1.0308758e-014             kt2=-0.042873075 lkt2=3.0723421e-009             wkt2=-2.5416844e-008            pkt2=4.4336207e-015 ute=-0.61639816                wute=-9.6263781e-008            ua1=3.411758e-009 lua1=-1.9592852e-016            wua1=-9.9993131e-016            pua1=-6.5479791e-023 ub1=-2.9256354e-18             lub1=7.1948561e-26              wub1=9.5903745e-25 pub1=1.2420305e-31              uc1=-5.6832829e-010            luc1=3.2198727e-017 wuc1=7.5154953e-016             puc1=-1.0238924e-022            at=162672.47 wat=-0.032535417               lcit=5.2229582e-010             wcit=5.1732994e-010 pcit=-2.1576837e-016            lu0=-1.9558933e-009            pu0=5.8042954e-016 lvsat=0.0017997505               pvsat=-5.2914334e-009            lpclm=9.042913e-008 ppclm=1.3711162e-014             lbigc=1.7841171e-010             pbigc=-1.6764482e-016 lbigsd=4.6070335e-013             pbigsd=-4.1490943e-018            lute=-4.5143609e-008 pute=5.0052259e-014             lat=-0.0032544114              pat=-7.0811685e-009 leta0=1.0169054e-010             peta0=-9.1582502e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00499996                 lvoff_mcl=2.66e-15                   wvoff_mcl=2e-15 pvoff_mcl=-5.7e-21                   u0_ff=-0.000726021               u0_ss=0.000454226 u0_fs=-0.000423829               u0_sf=0.000454226                wu0_ff=6.57775e-10 wu0_ss=-6.57775e-10               wu0_fs=3.83989e-10                wu0_sf=-6.57775e-10 pdiblc2_ff=-9.05987e-05               lpdiblc2_ff=4.04069e-11                wpdiblc2_ff=-4.7e-17 ppdiblc2_ff=2.9e-23                    lu0_ff=2.24629e-10                lu0_ss=-1.03409e-10 lu0_fs=8.98517e-11                lu0_sf=-1.03409e-10               pu0_ff=-2.03514e-16 pu0_ss=2.03514e-16                pu0_fs=-8.14057e-17               pu0_sf=2.03514e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.4 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.64340484 lvth0=-5.454483e-009             wvth0=-2.155959e-008             pvth0=6.8836022e-016 k2=-0.054305858               lk2=1.9033262e-009             wk2=-1.0261271e-008 pk2=-2.2095214e-015            cit=0.0045011297               voff=-0.19457119 lvoff=-2.0393825e-009            wvoff=-3.0957056e-008            pvoff=1.5547947e-015 eta0=0.041172395                weta0=-2.1893e-008               etab=-0.0072199256 wetab=-2.5187474e-009            u0=0.024039295                wu0=2.7100104e-009 ua=-1.1256042e-009            lua=-2.4569408e-017            wua=4.8169972e-017 pua=7.8107865e-024             ub=1.5445496e-018             lub=3.2090249e-027 wub=6.2052007e-026             pub=-3.4894986e-032            uc=6.24648e-011 luc=6.9888503e-018             wuc=-7.8065453e-017            puc=-1.2910334e-023 vsat=133050.32                  wvsat=-0.018716784               a0=1.8111491 la0=-3.9526599e-007            wa0=-6.1502224e-007            pa0=4.12487e-014 ags=1.2940506                  lags=8.0923927e-009             wags=1.8547807e-006 pags=-7.2880089e-014            keta=-0.13330724                lketa=-2.734725e-008 wketa=1.2487791e-008             pketa=2.0843705e-014             pclm=0.40707256 wpclm=9.2245598e-008             pdiblc2=0.001                      ppdiblc2=0 wpdiblc2=0                          lpdiblc2=0                          aigbacc=0.0088059516 laigbacc=-1.0496466e-010            waigbacc=-4.530101e-011             paigbacc=1.5163329e-018 aigc=0.0096482906               laigc=4.3212366e-011             waigc=-9.7380657e-011 paigc=-1.5748221e-018            bigc=0.0010525266               wbigc=-2.1452179e-010 aigsd=0.0096223733               laigsd=-2.2091765e-011            waigsd=-7.821935e-011 paigsd=1.8134481e-017             bigsd=0.00061530678              wbigsd=-8.5787084e-011 tvoff=0.000883933                ltvoff=1.02744e-010               wtvoff=2.88805e-010 ptvoff=-8.54126e-017              kt1=-0.19408089                lkt1=1.0550104e-008 wkt1=8.2785969e-008             pkt1=-8.3136926e-015            kt2=-0.02353809 lkt2=-1.0266747e-009            wkt2=-7.0785186e-009            pkt2=5.4589576e-016 ute=-0.94088649                wute=3.8002888e-007             ua1=4.3649176e-009 lua1=-3.9799836e-016            wua1=-2.4932071e-015            pua1=2.5109467e-022 ub1=-4.7353139e-18             lub1=4.556004e-25               wub1=3.1909718e-24 pub1=-3.4896701e-31             uc1=-7.5347107e-010            luc1=7.1448996e-017 wuc1=4.3549403e-016             puc1=-3.538547e-023             at=213495.92 wat=-0.11516804                lcit=-9.6590799e-012            wcit=-9.1077406e-010 pcit=8.6989674e-017             lu0=-3.1876396e-010            pu0=-2.9326948e-016 lvsat=-0.0018224043              pvsat=1.1917352e-009             lpclm=2.7849221e-008 ppclm=1.1475699e-014             lbigc=5.090799e-011              pbigc=-2.64992e-019 lbigsd=-7.4850369e-012            pbigsd=1.8186862e-017             lute=2.3647917e-008 pute=-5.0921784e-014            lat=-0.014028984               pat=1.0436947e-008 leta0=4.3462901e-011             peta0=5.8333223e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.005                      lvoff_mcl=2.56e-16                   wvoff_mcl=-3.6e-15 pvoff_mcl=-5.2e-22                   u0_ff=0.000356451                u0_ss=0.000163577 u0_sf=-5.64516e-05               u0_mc=7.62492e-05                wu0_ff=-5.08459e-10 wu0_ss=3.70951e-10                wu0_sf=5.08459e-10                wu0_mc=-6.87463e-10 pdiblc2_ff=0.000168254                ppdiblc2_ff=-3.7e-23                   wpdiblc2_ff=4.7e-16 lpdiblc2_ff=-1.44698e-11               lu0_ff=-4.85488e-12               lu0_ss=-4.17912e-11 lu0_sf=4.85484e-12                lu0_mc=-1.61648e-11               pu0_ff=4.37275e-17 pu0_ss=-1.45758e-17               pu0_sf=-4.37275e-17               pu0_mc=1.45742e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.5 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.57358496 lvth0=5.5002665e-010             wvth0=-1.8829797e-008            pvth0=4.5359813e-016 k2=-0.029306343               lk2=-2.4663199e-010            wk2=-4.6623718e-008 pk2=9.1764902e-016             cit=0.0034631975               voff=-0.20611269 lvoff=-1.0468131e-009            wvoff=-2.0997666e-008            pvoff=6.9828716e-016 eta0=0.042911317                weta0=-1.3710986e-008            etab=-0.0080909665 wetab=5.3283483e-009             u0=0.019656978                wu0=-1.5563369e-009 ua=-1.7916013e-009            lua=3.2706345e-017             wua=1.3411182e-016 pua=4.1978759e-025             ub=1.769823e-018              lub=-1.6164487e-026 wub=-2.9655465e-025            pub=-4.0548144e-033            uc=1.7843176e-010 luc=-2.984308e-018             wuc=-3.2599307e-016            puc=8.4114412e-024 vsat=100864.13                  wvsat=-0.014406721               a0=2.4709451 la0=-4.5200845e-007            wa0=9.6105397e-007             pa0=-9.4293854e-014 ags=1.3881482                  lags=0                          wags=1.0073378e-006 pags=0                          keta=-0.16881395                lketa=-2.4293673e-008 wketa=1.4992544e-007             pketa=9.0240676e-015             pclm=1.2665223 wpclm=-1.1068404e-008            pdiblc2=0.001                      aigbacc=0.0068245647 laigbacc=6.5434616e-011             waigbacc=-1.342535e-011             paigbacc=-1.2249739e-018 aigc=0.01039443                 laigc=-2.0955587e-011            waigc=-5.3487612e-010 paigc=3.6049788e-017             bigc=0.0018031095               wbigc=-7.5039803e-010 aigsd=0.0093154834               laigsd=4.3007642e-012             waigsd=2.5584226e-010 paigsd=-1.0594817e-017            bigsd=0.00051016578              wbigsd=2.515668e-010 tvoff=0.0019542                  ltvoff=1.07012e-011               wtvoff=-1.90344e-009 ptvoff=1.03121e-016               kt1=-0.12149994                lkt1=4.3081419e-009 wkt1=-5.4997705e-008            pkt1=3.5357033e-015             kt2=-0.053265024 lkt2=1.5298416e-009             wkt2=1.1614082e-008             pkt2=-1.0616679e-015 ute=-0.65625528                wute=-2.2083272e-007            ua1=2.0742457e-009 lua1=-2.0100058e-016            wua1=1.0382369e-015             pua1=-5.2609506e-023 ub1=-2.3154393e-018            lub1=2.4749119e-025             wub1=-1.666494e-024 pub1=6.8775047e-032             uc1=-2.5038778e-010            luc1=2.8183833e-017 wuc1=-2.6527681e-017            puc1=4.3483974e-024             at=77413.721 wat=0.01823829                 lcit=7.9603086e-011             wcit=-3.189903e-010 pcit=3.609627e-017              lu0=5.8115296e-011             pu0=7.3636392e-017 lvsat=0.00094560858              pvsat=8.2106983e-010             lpclm=-4.606346e-008 ppclm=2.0360703e-014             lbigc=-1.3642132e-011            pbigc=4.5820365e-017 lbigsd=1.5570886e-012             pbigsd=-1.0825572e-017            lute=-8.3036694e-010 pute=7.5231245e-016             lat=-0.0023259147              pat=-1.0359971e-009 leta0=-1.0608436e-010            peta0=-1.203209e-016             letab=7.4909514e-011 petab=-6.7485023e-016            jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499999 lvoff_mcl=2.56e-16                   wvoff_mcl=-3.5e-15                   pvoff_mcl=-1.2e-22 u0_ff=0.000716666                u0_ss=-0.0007701                 u0_mc=-0.000266872 wu0_ff=4.4e-16                    wu0_ss=4.81277e-10                wu0_mc=2.40612e-09 lu0_ff=-3.58334e-11               lu0_ss=3.85051e-11                lu0_mc=1.33436e-11 pu0_ff=-2.2e-23                   pu0_ss=-2.40639e-17               pu0_mc=-1.20306e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.6 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.54704882 lvth0=1.8768333e-009             wvth0=-2.5536974e-008            pvth0=7.8895694e-016 k2=-0.011595748               lk2=-1.1321617e-009            wk2=-6.50951e-008 pk2=1.8412182e-015             cit=0.0022709712               voff=-0.16501639 lvoff=-3.1016283e-009            wvoff=-6.8885171e-009            pvoff=-7.1702863e-018 eta0=0.026613416                weta0=-1.1528421e-008            etab=0.017228015 wetab=-1.755383e-008             u0=0.021878052                wu0=-5.3930627e-009 ua=-1.1697569e-009            lua=1.6141232e-018             wua=-7.0118818e-016 pua=4.2184788e-023             ub=1.3808556e-018             lub=3.283884e-027 wub=4.0256799e-025             pub=-3.9010946e-032            uc=5.2868061e-011 luc=3.2938768e-018             wuc=-2.8540699e-016            puc=6.3821374e-024 vsat=75963.579                  wvsat=0.027346005                a0=-2.4909972 la0=-2.0391134e-007            wa0=8.6290434e-006             pa0=-4.7769333e-013 ags=1.3881482                  lags=0                          wags=1.0073378e-006 pags=0                          keta=-1.2700367                 lketa=3.0767463e-008 wketa=8.0536655e-007             pketa=-2.3747988e-014            pclm=0.75522527 wpclm=3.6521591e-007             pdiblc2=0.001                      aigbacc=0.0086789935 laigbacc=-2.7286825e-011            waigbacc=-9.3977467e-011            paigbacc=2.802632e-018 aigc=0.011494975                laigc=-7.5982864e-011            waigc=7.0239177e-010 paigc=-2.5813607e-017            bigc=0.0032787953               wbigc=6.4096903e-010 aigsd=0.0083876165               laigsd=5.0694113e-011             waigsd=7.3985857e-010 paigsd=-3.4795632e-017            bigsd=-0.00033115422             wbigsd=7.5369013e-010 tvoff=0.00238967                 ltvoff=-1.10724e-011              wtvoff=-6.81144e-011 ptvoff=1.13544e-017               kt1=-0.10240762                lkt1=3.3535259e-009 wkt1=-4.0458407e-008            pkt1=2.8087384e-015             kt2=0.014953976 lkt2=-1.8811084e-009            wkt2=-1.4817832e-008            pkt2=2.5992779e-016 ute=-0.13711123                wute=-1.4249758e-006            ua1=1.1916178e-009 lua1=-1.5686918e-016            wua1=1.3155342e-017             pua1=-1.3554296e-024 ub1=5.1217018e-019             lub1=1.0611071e-025             wub1=-2.3206014e-024 pub1=1.0148041e-031             uc1=-4.5953077e-011            luc1=1.7962098e-017 wuc1=1.3586748e-017             puc1=2.3426759e-024             at=13524.794 wat=0.042009451                lcit=1.392144e-010              wcit=8.6183343e-010 pcit=-2.2944916e-017            lu0=-5.2938424e-011            pu0=2.6547268e-016 lvsat=0.0021906359               pvsat=-1.2665665e-009            lpclm=-2.0498606e-008 ppclm=1.5464873e-015             lbigc=-8.7426426e-011            pbigc=-2.3747988e-017 lbigsd=4.3623089e-011             pbigsd=-3.5931739e-017            lute=-2.678757e-008 pute=6.0959468e-014             lat=0.00086853168              pat=-2.2245552e-009 leta0=7.088107e-010              peta0=-2.2944916e-016            letab=-1.1910396e-009 petab=4.6925866e-016             jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499997 lvoff_mcl=-1.76e-15                  wvoff_mcl=3e-14                      pvoff_mcl=-6.5e-21 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.7 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.58787066 lvth0=2.0313774e-010             wvth0=-2.6409753e-008            pvth0=8.2474087e-016 k2=0.026573387                lk2=-2.6970963e-009            wk2=-5.6488061e-008 pk2=1.4883295e-015             cit=0.00076583539              voff=-0.17234528 lvoff=-2.8011438e-009            wvoff=-2.0359401e-008            pvoff=5.4513596e-016 eta0=0.029305268                weta0=-4.5777906e-008            etab=-0.0052783334 wetab=-3.8716793e-008            u0=0.029796553                wu0=-5.9059095e-009 ua=-7.9929337e-010            lua=-1.3574881e-017            wua=-1.0486948e-015 pua=5.6432557e-023             ub=1.4479625e-018             lub=5.3250069e-028 wub=4.1021089e-025             pub=-3.9324305e-032            uc=3.5493996e-010 luc=-9.0910713e-018            wuc=-2.1012287e-016            puc=3.2954883e-024 vsat=113584.55                  wvsat=-0.053296459               a0=14.030274 la0=-8.8128347e-007            wa0=-2.0486116e-005            pa0=7.1602823e-013 ags=1.3881482                  lags=0                          wags=1.0073378e-006 pags=0                          keta=-0.38746128                lketa=-5.4181281e-009 wketa=4.9297992e-007             pketa=-1.0940136e-014            pclm=0.75586226 wpclm=6.9770453e-007             pdiblc2=0.001                      aigbacc=0.0079934338 laigbacc=8.2112437e-013             waigbacc=-1.6923393e-010            paigbacc=5.8881471e-018 aigc=0.0099094043               laigc=-1.0974462e-011            waigc=9.0311523e-010 paigc=-3.4043268e-017            bigc=0.0014159456               wbigc=9.8724698e-010 aigsd=0.010029982                laigsd=-1.6642883e-011            waigsd=-1.1815724e-009 paigsd=4.3983035e-017             bigsd=0.0012783577               wbigsd=-1.2956826e-009 tvoff=0.000893781                ltvoff=5.02591e-011               wtvoff=2.18983e-009 ptvoff=-8.12213e-017              kt1=-0.16189465                lkt1=5.7924941e-009 wkt1=1.1550076e-007             pkt1=-3.5855875e-015            kt2=-0.076948306 lkt2=1.8868852e-009             wkt2=-2.9396623e-008            pkt2=8.5765822e-016 ute=-0.31153296                wute=-5.2415254e-007            ua1=-1.7871252e-009 lua1=-3.474072e-017             wua1=1.3429294e-016             pua1=-6.3220711e-024 ub1=1.9981757e-018             lub1=4.5184484e-026             wub1=2.0850264e-025 pub1=-2.2128503e-033            uc1=9.7977616e-010             luc1=-2.40928e-017 wuc1=1.7557157e-016             puc1=-4.2987016e-024            at=72578.801 wat=-0.058832612               lcit=2.0092497e-010             wcit=2.8093531e-009 pcit=-1.0279322e-016            lu0=-3.7759695e-010            pu0=2.864994e-016 lvsat=0.00064817604              pvsat=2.0397746e-009             lpclm=-2.0524723e-008 ppclm=-1.2085546e-014            lbigc=-1.1049588e-011            pbigc=-3.7945384e-017 lbigsd=-2.23669e-011              pbigsd=4.8092544e-017             lute=-1.9636278e-008 pute=2.4025713e-014             lat=-0.0015526826              pat=1.9099694e-009 leta0=5.9844477e-010             peta0=1.1747797e-015             letab=-2.6827928e-010 petab=1.3369402e-015             jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_ff=-0.00987137 voff_ss=0.0177778                  voff_mcl=-0.0029055                 voff_mc='-0.0197638+0.00198603' lvoff_ff=4.04726e-10                lvoff_ss=-7.28888e-10               lvoff_mcl=3.24126e-10 lvoff_mc='8.10316e-10-8.1427e-11'   wvoff_ff=-7.16321e-09               wvoff_ss=5e-15 wvoff_mcl=7.16239e-09                wvoff_mc='1.7906e-08-1.7906e-08'    pvoff_ff=2.93691e-16 pvoff_ss=-2e-22                     pvoff_mcl=-2.93664e-16               pvoff_mc='-7.34146e-16+7.34146e-16' u0_mc=0.000397205                wu0_mc=-3.5812e-09                ua_ff=7.95293e-12 ua_ss=-7.95293e-12               lua_ff=-3.2607e-19                lua_ss=3.2607e-19 wua_ff=-7.1632e-17                wua_ss=7.1632e-17                 pua_ff=2.93691e-24 pua_ss=-2.93691e-24               vsat_ff=-795.293                   vsat_ss=397.646 wvsat_ff=0.0071632                  wvsat_ss=-0.0035816                 ua1_fs=-7.9064e-11 ua1_sf=7.9064e-11                 lua1_fs=3.24163e-18                lua1_sf=-3.24163e-18 wua1_fs=7.1632e-17                 wua1_sf=-7.1632e-17                pua1_fs=-2.93691e-24 pua1_sf=2.93691e-24                lu0_mc=-1.62854e-11               pu0_mc=1.46829e-16 lvsat_ff=3.2607e-05                 lvsat_ss=-1.63035e-05               pvsat_ff=-2.93691e-10 pvsat_ss=1.46846e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_hvt_mac.8 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=0.6169285 lvth0=2.9787052e-012             wvth0=-1.5980844e-008            pvth0=5.4695396e-019 k2=-0.049797261               lk2=1.1494897e-009             wk2=1.9655439e-010 pk2=-1.7805647e-015            cit=0.0039546517               voff=-0.23559317 lvoff=0                          wvoff=1.5513589e-008             pvoff=0 eta0=0.0163484                  weta0=5.5733496e-009             etab=0.0051666667 wetab=-1.3741e-008               u0=0.025731517                wu0=3.5438039e-009 ua=-1.3243532e-009            lua=1.5742588e-016             wua=2.2188744e-016 pua=-9.3108273e-024            ub=1.8606003e-018             lub=-6.8870118e-030 wub=6.224255e-027              pub=3.7603085e-036             uc=6.509409e-010 luc=-4.4926837e-016            wuc=-8.9358592e-017            puc=6.2185677e-023 vsat=147750                     wvsat=-0.0206115                 a0=-0.035655305 la0=-1.5253093e-011            wa0=4.7546492e-007             pa0=1.0501516e-017 ags=-0.45556576                lags=3.2442921e-006             wags=1.0252632e-006 pags=-9.8482483e-013            keta=0.088539367                lketa=-2.5882994e-007 wketa=-3.7309496e-008            pketa=5.805318e-014              pclm=0.4 wpclm=0                          pdiblc2=0.0010037276               lpdiblc2=-3.3533238e-011 wpdiblc2=-8.074958e-012             ppdiblc2=7.2642322e-017             aigbacc=0.010732764 laigbacc=-1.3878893e-009            waigbacc=1.5950396e-011             paigbacc=-2.5858342e-018 aigc=0.010542695                laigc=2.0918639e-010             waigc=-4.3648974e-010 paigc=-1.1873915e-016            bigc=0.0021989383               wbigc=-6.3387233e-010 aigsd=0.0094741356               laigsd=5.5114053e-011             waigsd=1.6665244e-011 paigsd=-4.6438278e-017            bigsd=0.00059131242              wbigsd=-6.1765795e-012 tvoff=0.0015506                  ltvoff=-3.30749e-010              wtvoff=2.61182e-010 ptvoff=3.49219e-017               kt1=-0.10632645                lkt1=-1.246545e-011 wkt1=-2.2405734e-009            pkt1=7.1104014e-018             kt2=-0.018504655 lkt2=4.9585158e-013             wkt2=-1.0091342e-008            pkt2=-4.3373449e-019 ute=-0.675                     ua1=1.0497307e-009             lua1=-1.0881562e-020 wua1=9.7743778e-016             pua1=6.9736629e-027             ub1=-8.347e-020 wub1=-1.2803864e-024            uc1=4.6540998e-011             luc1=-5.5381578e-016 wuc1=-9.2483657e-017            puc1=3.0238337e-022             at=75106.517 wat=0.040891842                lcit=0                          wcit=4.108559e-011 pcit=0                          lu0=0                          pu0=0 lvsat=0                          pvsat=0                          lpclm=0 ppclm=0                          lat=0                          pat=0 leta0=0                          peta0=0                          jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00166855 voff_mc=0.00139022                 lvoff_mcl=2.98495e-09                lvoff_mc=-1.25203e-08 wvoff_mcl=5.06e-15                   wvoff_mc=-7.59059e-10               pvoff_mcl=4.8e-21 pvoff_mc=6.83608e-15 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.9 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.61627502 lvth0=5.8850176e-010             wvth0=-1.7075135e-008            pvth0=9.8103191e-016 k2=-0.038263057               lk2=-9.1851575e-009            wk2=-5.4335627e-009 pk2=3.2640202e-015             cit=0.0047025953               voff=-0.2445037 lvoff=7.9838422e-009             wvoff=2.3068242e-008             pvoff=-6.7689689e-015 eta0=0.0163484                  weta0=5.5733496e-009             etab=0.0051666667 wetab=-1.3741e-008               u0=0.023715002                wu0=7.5150628e-009 ua=-1.4092387e-009            lua=2.3348324e-016             wua=5.2973638e-016 pua=-2.8514347e-022            ub=1.9419108e-018             lub=-7.2861168e-026 wub=3.6506918e-026             pub=-2.7129506e-032            uc=2.0489525e-010 luc=-4.9611462e-017            wuc=-3.2341085e-017            puc=1.1097991e-023 vsat=160221.48                  wvsat=-0.027420929               a0=-0.29654872 la0=2.3374525e-007             wa0=7.1750237e-007             pa0=-2.1685506e-013 ags=3.6297597                  lags=-4.1615951e-007            wags=-4.1946375e-007 pags=3.0965055e-013             keta=-0.28015792                lketa=7.1522828e-008 wketa=6.3885207e-008             pketa=-3.2617273e-014            pclm=0.45366454 wpclm=-8.3415504e-008            pdiblc2=0.00089194934              lpdiblc2=6.6620057e-011 wpdiblc2=-5.3077513e-011            ppdiblc2=1.1296461e-016             aigbacc=0.0096198358 laigbacc=-3.9070528e-010            waigbacc=1.1258492e-011             paigbacc=1.6181121e-018 aigc=0.012103561                laigc=-1.1893498e-009            waigc=-1.408234e-009 paigc=7.5194374e-016             bigc=0.0036637345               wbigc=-1.5762973e-009 aigsd=0.0094558605               laigsd=7.1488526e-011             waigsd=1.7982099e-011 paigsd=-4.7618181e-017            bigsd=0.0004986324               wbigsd=7.2674564e-011 tvoff=0.000423906                ltvoff=6.78769e-010               wtvoff=7.70369e-010 ptvoff=-4.2131e-016               kt1=-0.13173841                lkt1=2.275665e-008 wkt1=1.3025483e-008             pkt1=-1.3671276e-014            kt2=0.012540583 lkt2=-2.7816038e-008            wkt2=-1.7185617e-008            pkt2=6.3560363e-015 ute=-0.65222146                wute=1.8113081e-009             ua1=1.1000357e-009 lua1=-4.5084125e-017            wua1=1.3106531e-015             pua1=-2.9855397e-022 ub1=3.0042367e-019             lub1=-3.4396873e-025            wub1=-1.7164622e-024 pub1=3.9072394e-031             uc1=-1.1596351e-009            luc1=5.2691798e-016 wuc1=4.3555314e-016             puc1=-1.7073761e-022            at=67206.113 wat=0.064482772                lcit=-6.7015751e-010            wcit=8.1805975e-011 pcit=-3.6485465e-017            lu0=1.8067971e-009             pu0=-3.558248e-015 lvsat=-0.011174447               pvsat=6.1012483e-009             lpclm=-4.8083425e-008 ppclm=7.4740291e-014             lbigc=-1.3124574e-009            pbigc=8.4441276e-016 lbigsd=8.3041293e-011             pbigsd=-7.0650625e-017            lute=-2.0409573e-008 pute=-1.622932e-015             lat=0.007078762                pat=-2.1137473e-008 leta0=0                          peta0=0                          jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499997 voff_mc=-0.0250548                 lvoff_mcl=5.04e-14                   lvoff_mc=1.11744e-08 wvoff_mcl=3.11e-14                   wvoff_mc=1.36799e-08                pvoff_mcl=-1.7e-21 pvoff_mc=-6.10125e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.10 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.61764568 lvth0=-2.2812973e-011            wvth0=-1.1874893e-008            pvth0=-1.3382762e-015 k2=-0.046683195               lk2=-5.4297756e-009            wk2=1.9603314e-010 pk2=7.5322045e-016             cit=0.0024211084               voff=-0.21040285 lvoff=-7.2251369e-009            wvoff=3.3694651e-009             pvoff=2.0166855e-015 eta0=0.021478528                weta0=2.7722996e-009             etab=0.0051666667 wetab=-1.3741e-008               u0=0.028493213                wu0=1.5499496e-009 ua=-7.8608188e-010            lua=-4.4444693e-017            wua=-8.4180121e-017 pua=-1.1336716e-023            ub=2.0336154e-018             lub=-1.1376141e-025 wub=-4.9009567e-027            pub=-8.6615935e-033            uc=2.4757661e-010 luc=-6.8647349e-017            wuc=-2.9220189e-017            puc=9.706071e-024 vsat=166211.68                  wvsat=-0.033659578               a0=1.4072602 la0=-5.2615355e-007            wa0=-1.6550646e-008            pa0=1.1053259e-013 ags=2.4218518                  lags=1.2256741e-007             wags=5.2380222e-007 pags=-1.1104607e-013            keta=-0.060263264               lketa=-2.6550188e-008 wketa=-5.4973278e-008            pketa=2.0393611e-014             pclm=-0.002477386 wpclm=1.8531265e-007             pdiblc2=0.0024528325               lpdiblc2=-6.2953382e-010 wpdiblc2=-8.6332119e-010            ppdiblc2=4.7433329e-016             aigbacc=0.0091787851 laigbacc=-1.9399664e-010            waigbacc=2.4251178e-011             paigbacc=-4.176626e-018 aigc=0.0098557227               laigc=-1.8681381e-010            waigc=-9.6029613e-011 paigc=1.6670057e-016             bigc=0.0012338276               wbigc=-1.3415092e-010 aigsd=0.0096006306               laigsd=6.921049e-012              waigsd=-8.1370518e-011 paigsd=-3.3069131e-018            bigsd=0.00077979207              wbigsd=-1.6340927e-010 tvoff=0.00254857                 ltvoff=-2.6883e-010               wtvoff=-3.01093e-010 ptvoff=5.65625e-017               kt1=-0.10786333                lkt1=1.2108364e-008 wkt1=3.7304295e-009             pkt1=-9.5256821e-015            kt2=-0.073195259 lkt2=1.0422148e-008             wkt2=2.0550552e-009             pkt2=-2.2253034e-015 ute=-1.0497094                 wute=2.9631621e-007             ua1=1.8857227e-009 lua1=-3.9550055e-016            wua1=3.8265661e-016             pua1=1.1533247e-022 ub1=-1.7436557e-018            lub1=5.6769067e-025             wub1=-1.1183613e-025 pub1=-3.2493929e-031            uc1=1.2723048e-010             luc1=-4.7024059e-017 wuc1=1.2137329e-016             puc1=-3.0613392e-023            at=132659.13 wat=-0.005343336               lcit=3.4738566e-010             wcit=1.2847483e-010 pcit=-5.7299773e-017            lu0=-3.2428508e-010            pu0=-8.9780748e-016 lvsat=-0.013846076               pvsat=8.8836857e-009             lpclm=1.5535587e-007 ppclm=-4.5112466e-014            lbigc=-2.2871886e-010            pbigc=2.0121548e-016 lbigsd=-4.2355919e-011            pbigsd=3.4642765e-017             lute=1.5687005e-007 pute=-1.3297212e-013            lat=-0.022113285               pat=1.0004971e-008 leta0=-2.2880372e-009            peta0=1.2492683e-015 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00499997                 lvoff_mcl=-5.2e-15                   wvoff_mcl=-3.56e-14 pvoff_mcl=1.8e-21                    u0_ff=0.000412222                u0_ss=-0.000684017 u0_fs=0.000274815                u0_sf=-0.000684017               wu0_ff=-3.73473e-10 wu0_ss=3.73473e-10                wu0_fs=-2.48982e-10               wu0_sf=3.73473e-10 pdiblc2_ff=-0.000228006               lpdiblc2_ff=1.01691e-10                wpdiblc2_ff=1.24491e-10 ppdiblc2_ff=-5.5523e-17                lu0_ff=-1.83851e-10               lu0_ss=3.05072e-10 lu0_fs=-1.22567e-10               lu0_sf=3.05072e-10                pu0_ff=1.66569e-16 pu0_ss=-1.66569e-16               pu0_fs=1.11046e-16                pu0_sf=-1.66569e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.11 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.64843605 lvth0=-6.5503723e-009            wvth0=-2.6117874e-008            pvth0=1.6812359e-015 k2=-0.06797038                lk2=-9.1689257e-010            wk2=2.118786e-009 pk2=3.4559684e-016             cit=0.0032416188               voff=-0.25060432 lvoff=1.2975735e-009             wvoff=1.980896e-008              pvoff=-1.4684875e-015 eta0=0.00091595873              weta0=1.4579332e-008             etab=0.0051666667 wetab=-1.3741e-008               u0=0.032497121                wu0=-4.9527799e-009 ua=-8.3131895e-010            lua=-3.4854435e-017            wua=-2.1845246e-016 pua=1.7129021e-023             ub=1.673586e-018              lub=-3.7435167e-026 wub=-5.4854944e-026            pub=1.9286519e-033             uc=-2.5805816e-011 luc=-1.0690275e-017            wuc=1.9077258e-018             puc=3.1069531e-024 vsat=98637.427                  wvsat=0.012461299                a0=-0.70126247 la0=-7.9146734e-008            wa0=1.6612226e-006             pa0=-2.4515535e-013 ags=3.8588624                  lags=-1.8207884e-007            wags=-4.6893889e-007 pags=9.9415044e-014             keta=-0.20487844                lketa=4.1082291e-009 wketa=7.7331294e-008             pketa=-7.6549584e-015            pclm=0.53454318 wpclm=-2.3242792e-008            pdiblc2=-0.00051666667             ppdiblc2=0 lpdiblc2=0                          wpdiblc2=1.3741e-009                aigbacc=0.0087890962 laigbacc=-1.113826e-010             waigbacc=-3.0030032e-011            paigbacc=7.3309906e-018 aigc=0.008311837                laigc=1.4048995e-010             waigc=1.1134463e-009 paigc=-8.9708317e-017            bigc=-0.00065055127             wbigc=1.3284668e-009 aigsd=0.0095301756               laigsd=2.1857517e-011             waigsd=5.311818e-012 paigsd=-2.1683568e-017            bigsd=0.00044857016              wbigsd=6.5276293e-011 tvoff=0.00149411                 ltvoff=-4.52847e-011              wtvoff=-2.64013e-010 ptvoff=4.87014e-017               kt1=0.00039096149              lkt1=-1.0841545e-008 wkt1=-9.3405529e-008            pkt1=1.1067141e-014             kt2=-0.013885969 lkt2=-2.1514215e-009            wkt2=-1.582334e-008             pkt2=1.5649163e-015 ute=0.28876874                 wute=-7.3403877e-007            ua1=-8.1524545e-010 lua1=1.771047e-016              wua1=2.2000206e-015             pua1=-2.699487e-022 ub1=3.0755886e-018             lub1=-4.5398913e-025            wub1=-3.8857059e-024 pub1=4.7512111e-031             uc1=-8.9094951e-011            luc1=-1.1630682e-018 wuc1=-1.6643073e-016            puc1=3.0401061e-023             at=-14085.759 wat=0.091020966                lcit=1.7343745e-010             wcit=2.3034278e-010 pcit=-7.8895779e-017            lu0=-1.1731134e-009            pu0=4.8077116e-016 lvsat=0.00047966559              pvsat=-8.9394008e-010            lpclm=4.1507511e-008 ppclm=-8.98712e-016              lbigc=1.7076945e-010             pbigc=-1.0885947e-016 lbigsd=2.7863126e-011             pbigsd=-1.3838574e-017            lute=-1.2688732e-007 pute=8.5463137e-014             lat=0.0089966322               pat=-1.0424261e-008 leta0=2.0712276e-009             peta0=-1.2538225e-015 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00500007                 lvoff_mcl=-6.3e-15                   wvoff_mcl=-8.9e-15 pvoff_mcl=-5.6e-22                   u0_ff=-0.000970314               u0_ss=0.00144209 u0_fs=-0.00051037                u0_sf=0.00127032                 u0_mc=-0.00171772 wu0_ff=6.93593e-10                wu0_ss=-7.87381e-10               wu0_fs=4.62396e-10 wu0_sf=-6.93593e-10               wu0_mc=9.37878e-10                pdiblc2_ff=0.000423439 ppdiblc2_ff=1.9883e-17                 lpdiblc2_ff=-3.64158e-11               wpdiblc2_ff=-2.31198e-10 lu0_ff=1.09247e-10                lu0_ss=-1.45663e-10               lu0_fs=4.38919e-11 lu0_sf=-1.09247e-10               lu0_mc=3.64158e-10                pu0_ff=-5.9649e-17 pu0_ss=7.9532e-17                 pu0_fs=-3.9766e-17                pu0_sf=5.9649e-17 pu0_mc=-1.9883e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.12 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.55369095 lvth0=1.5977064e-009             wvth0=-8.058334e-010             pvth0=-4.9559964e-016 k2=-0.09921774                lk2=1.7703804e-009             wk2=1.6716008e-008 pk2=-9.0976422e-016            cit=0.0036339398               voff=-0.23469938 lvoff=-7.0251111e-011            wvoff=4.9018735e-009             pvoff=-1.86478e-016 eta0=0.040416667                weta0=-1.1450833e-008            etab=0.029315716 wetab=-2.8562106e-008            u0=0.015996822                wu0=1.7597641e-009 ua=-1.3207596e-009            lua=7.2374564e-018             wua=-2.9247083e-016 pua=2.34946e-023               ub=1.0574183e-018             lub=1.555525e-026 wub=3.4888399e-025             pub=-3.2792897e-032            uc=-4.3153836e-010 luc=2.4202724e-017             wuc=2.2663985e-016             puc=-1.622001e-023 vsat=83726.415                  wvsat=0.0011200442               a0=7.2113804 la0=-7.5963402e-007            wa0=-3.3337803e-006            pa0=1.8441491e-013 ags=1.7416667                  lags=0                          wags=6.8705e-007 pags=0                          keta=0.0759125                  lketa=-2.0039792e-008 wketa=-7.1796725e-008            pketa=5.1700512e-015             pclm=1.0851012 wpclm=1.5329918e-007             pdiblc2=-0.00051666667             wpdiblc2=1.3741e-009 aigbacc=0.0063416641               laigbacc=9.9096559e-011             waigbacc=4.2408258e-010 paigbacc=-3.1722694e-017            aigc=0.0095382905               laigc=3.5014956e-011 waigc=2.4078589e-010             paigc=-1.4659524e-017            bigc=0.00067082287 wbigc=2.7545361e-010             aigsd=0.01004524                 laigsd=-2.2438026e-011 waigsd=-4.0531719e-010            paigsd=1.3630527e-017             bigsd=0.00091782852 wbigsd=-1.1777564e-010            tvoff=-0.00127859                ltvoff=1.93167e-010 wtvoff=1.02546e-009               ptvoff=-6.21931e-017              kt1=-0.29987363 lkt1=1.498121e-008              wkt1=1.0660886e-007             pkt1=-6.1340965e-015 kt2=-0.051440455               lkt2=1.0782643e-009             wkt2=9.9610223e-009 pkt2=-6.5253881e-016            ute=-1.1108529                 wute=1.9103273e-007 ua1=7.5362726e-009             lua1=-5.4112585e-016            wua1=-3.9103595e-015 pua1=2.5554399e-022             ub1=-1.0210403e-017            lub1=6.8860615e-025 wub1=5.4863431e-024             pub1=-3.3087511e-031            uc1=-7.0501859e-010 luc1=5.1806364e-017             wuc1=3.8536783e-016             puc1=-1.7053616e-023 at=194235.86                  wat=-0.087602566               lcit=1.3969784e-010 wcit=-4.7368281e-010            pcit=-1.8349579e-017            lu0=2.4591223e-010 pu0=-9.6507619e-017            lvsat=0.0017620126               pvsat=8.1407791e-011 lpclm=-5.840475e-009             ppclm=-1.6081321e-014            lbigc=5.7131273e-011 pbigc=-1.830034e-017             lbigsd=-1.2493093e-011            pbigsd=1.9038919e-018 lute=-6.5198551e-009            pute=5.9069887e-015             lat=-0.0089190269 pat=4.9373626e-009             leta0=-1.3258333e-009            peta0=9.8477167e-016 letab=-2.0768182e-009            petab=1.2746151e-015 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00499997                 lvoff_mcl=-1.04e-15                  wvoff_mcl=-4.11e-14 pvoff_mcl=6e-23                      u0_ff=0.000716666                u0_ss=-0.000601204 u0_mc=0.00601204                 wu0_ff=-3.3e-16                   wu0_ss=3.28257e-10 wu0_mc=-3.28257e-09               lu0_ff=-3.58334e-11               lu0_ss=3.00602e-11 lu0_mc=-3.00602e-10               pu0_ff=1.7e-23                    pu0_ss=-1.64129e-17 pu0_mc=1.64129e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.13 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.5065664 lvth0=3.9539339e-009             wvth0=1.1140099e-008             pvth0=-1.0928962e-015 k2=-0.09487826                lk2=1.5534064e-009             wk2=1.0358855e-008 pk2=-5.9190658e-016            cit=-0.00090868045             voff=-0.16814709 lvoff=-3.3978659e-009            wvoff=-4.0521064e-009            pvoff=2.6122099e-016 eta0=0.014181502                weta0=-2.6510725e-010            etab=0.025237413 wetab=-2.4810344e-008            u0=0.011608675                wu0=3.910994e-009 ua=-2.3616349e-009            lua=5.9281223e-017             wua=3.7865329e-016 pua=-1.0061605e-023            ub=2.3460527e-018             lub=-4.8876468e-026 wub=-4.719006e-025             pub=8.2463329e-033             uc=-8.1511574e-012 luc=3.0333641e-018             wuc=-2.3012358e-016            puc=6.6181618e-024 vsat=199014.21                  wvsat=-0.084137864               a0=24.904035 la0=-1.6442667e-006            wa0=-1.6190855e-005            pa0=8.2726866e-013 ags=1.7416667                  lags=0                          wags=6.8705e-007 pags=0                          keta=-0.17879957                lketa=-7.304188e-009 wketa=-1.8329425e-007            pketa=1.0744928e-014             pclm=0.86296419 wpclm=2.6760445e-007             pdiblc2=-0.00051666667             wpdiblc2=1.3741e-009 aigbacc=0.0087710662               laigbacc=-2.2373544e-011            waigbacc=-1.773953e-010 paigbacc=-1.6488002e-018            aigc=0.014376885                laigc=-2.0691474e-010 waigc=-1.9086181e-009            paigc=9.2810676e-017             bigc=0.0065109332 wbigc=-2.2873479e-009            aigsd=0.0094430677               laigsd=7.6705896e-012 waigsd=-2.1638026e-010            paigsd=4.1836798e-018             bigsd=0.00082109492 wbigsd=-2.902476e-010             tvoff=0.00449114                 ltvoff=-9.53191e-011 wtvoff=-1.97204e-009              ptvoff=8.76819e-017               kt1=0.038525394 lkt1=-1.9387411e-009            wkt1=-1.6814372e-007            pkt1=7.6035324e-015 kt2=0.024964243                lkt2=-2.7419706e-009            wkt2=-2.3887134e-008 pkt2=1.039869e-015              ute=-3.2795794                 wute=1.4221004e-006 ua1=-7.8619583e-009            lua1=2.287857e-016              wua1=8.2156953e-015 pua1=-3.5075875e-022            ub1=8.0528448e-018             lub1=-2.2455624e-025 wub1=-9.1524526e-024            pub1=4.0106467e-031             uc1=6.9705665e-010 luc1=-1.8297397e-017            wuc1=-6.5958006e-016            puc1=3.5193779e-023 at=-47400.341                 wat=0.097207623                lcit=3.6682886e-010 wcit=3.7425978e-009             pcit=-2.2916361e-016            lu0=4.6531962e-010 pu0=-2.0406912e-016            lvsat=-0.004002377               pvsat=4.3443032e-009 lpclm=5.2663741e-009             ppclm=-2.1796585e-014            lbigc=-2.3487424e-010 pbigc=1.0983973e-016             lbigsd=-7.6564126e-012            pbigsd=1.052749e-017 lute=1.0191647e-007             pute=-5.5646393e-014            lat=0.003162783 pat=-4.3031469e-009            leta0=-1.4075087e-011            peta0=4.2548536e-016 letab=-1.8729031e-009            petab=1.087027e-015 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.005                      lvoff_mcl=5.2e-15                    wvoff_mcl=5.6e-14 pvoff_mcl=7.2e-21                    ua1_fs=1.38185e-10                lua1_fs=-6.90926e-18 wua1_fs=-1.25196e-16               pua1_fs=6.25979e-24 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.14 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.65029918 lvth0=-1.9391099e-009            wvth0=-8.2969985e-008            pvth0=2.7656172e-015 k2=-0.014599911               lk2=-1.7380059e-009            wk2=-1.9185053e-008 pk2=6.1939365e-016             cit=0.013152551                voff=-0.18744718 lvoff=-2.6065619e-009            wvoff=-6.6770771e-009            pvoff=3.6884479e-016 eta0=-0.055892613               weta0=3.1411374e-008             etab=-0.06590336 wetab=1.620948e-008              u0=0.035574349                wu0=-1.1140592e-008 ua=-2.5273633e-009            lua=6.6076087e-017             wua=5.1693657e-016 pua=-1.573122e-023             ub=2.6102066e-018             lub=-5.9706779e-026 wub=-6.427823e-025             pub=1.5252483e-032             uc=4.0334116e-010 luc=-1.3837821e-017            wuc=-2.5397435e-016            puc=7.5960435e-024 vsat=45587.31                   wvsat=0.0083090409               a0=-17.891968 la0=1.1036938e-007             wa0=8.435435e-006              pa0=-1.8240925e-013 ags=1.7416667                  lags=0                          wags=6.8705e-007 pags=0                          keta=0.16176772                 lketa=-2.1267447e-008 wketa=-4.6215563e-009            pketa=3.4193471e-015             pclm=2.0570147 wpclm=-4.8113959e-007            pdiblc2=-0.00051666667             wpdiblc2=1.3741e-009 aigbacc=0.0083976414               laigbacc=-7.0631304e-012            waigbacc=-5.3544608e-010 paigbacc=1.3031282e-017             aigc=0.008810158                laigc=2.1321045e-011 waigc=1.8990324e-009             paigc=-6.3302997e-017            bigc=0.00038684942 wbigc=1.9196082e-009             aigsd=0.0085366028               laigsd=4.4835652e-011 waigsd=1.7142944e-010             paigsd=-1.1716518e-017            bigsd=-0.00058792307 wbigsd=3.9516777e-010             tvoff=0.00433062                 ltvoff=-8.87378e-011 wtvoff=-9.23945e-010              ptvoff=4.47099e-017               kt1=-0.056278838 lkt1=1.9482324e-009             wkt1=1.9812839e-008             pkt1=-1.0268636e-016 kt2=-0.15645845                lkt2=4.6963599e-009             wkt2=4.263957e-008 pkt2=-1.6877259e-015            ute=-1.9048341                 wute=9.1937825e-007 ua1=-2.2899075e-009            lua1=3.3161174e-019             wua1=5.8981375e-016 pua1=-3.8097604e-023            ub1=1.3759107e-018             lub1=4.9198056e-026 wub1=7.7227474e-025             pub1=-5.8491467e-033            uc1=8.0484116e-010 luc1=-2.2716562e-017            wuc1=3.3406267e-016             puc1=-5.5455732e-024 at=25026.191                  wat=-0.015749947               lcit=-2.0968163e-010 wcit=-8.413011e-009             pcit=2.6921635e-016             lu0=-5.1727302e-010 pu0=4.1304591e-016             lvsat=0.0022881258               pvsat=5.539801e-010 lpclm=-4.3689697e-008            ppclm=8.9019206e-015             lbigc=1.6213192e-011 pbigc=-6.2645463e-017            lbigsd=5.0113325e-011             pbigsd=-1.757454e-017 lute=4.5551911e-008             pute=-3.5034787e-014            lat=0.00019329523 pat=3.2811349e-010             leta0=2.8589636e-009             peta0=-8.7325037e-016 letab=1.8638686e-009             petab=-5.9478579e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_ff=-0.0339555                 voff_ss=0.0339555                  voff_mcl=0.00500006 voff_mc=-0.0447407                 lvoff_ff=1.39218e-09                lvoff_ss=-1.39218e-09 lvoff_mcl=-1.5e-15                   lvoff_mc=1.83437e-09                wvoff_ff=1.4657e-08 wvoff_ss=-1.4657e-08                wvoff_mcl=5.6e-14                    wvoff_mc=2.44284e-08 pvoff_ff=-6.00944e-16               pvoff_ss=6.00944e-16                pvoff_mcl=6.2e-21 pvoff_mc=-1.00157e-15               u0_mc=-0.00355556                wu0_mc=1.1e-15 ua_ff=-1.25037e-10               ua_ss=1.78963e-10                lua_ff=5.12652e-18 lua_ss=-7.33748e-18               wua_ff=4.88569e-17                wua_ss=-9.77138e-17 pua_ff=-2.00313e-24               pua_ss=4.00626e-24                vsat_ff=9807.41 vsat_ss=-8948.15                   vsat_fs=5392.59                    vsat_mc=-21570.4 wvsat_ff=-0.00244285                wvsat_ss=0.00488569                 wvsat_fs=-0.00488569 wvsat_mc=0.0195428                  ua1_fs=-1.38185e-10               lua1_fs=4.42193e-18 wua1_fs=1.25196e-16                pua1_fs=-4.00626e-24               lu0_mc=1.45778e-10 pu0_mc=2.4e-22                    lvsat_ff=-0.000402104               lvsat_ss=0.000366874 lvsat_fs=-0.000221096               lvsat_mc=0.000884385                pvsat_ff=1.00156e-10 pvsat_ss=-2.00313e-10               pvsat_fs=2.00313e-10                pvsat_mc=-8.01253e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.15 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.60591791 lvth0=-1.3986966e-008            wvth0=-9.9690601e-009            pvth0=7.6390567e-015 k2=-0.051043158               lk2=-2.608421e-009             wk2=8.7681387e-010 pk2=2.7125452e-016             cit=0.0049137437               voff=-0.22083871 lvoff=8.3846346e-009             wvoff=7.457654e-009              pvoff=-4.5780105e-015 eta0=0.022963911                weta0=1.9612805e-009             etab=-0.0128608 wetab=-3.8980032e-009            u0=0.032935248                wu0=-3.8943313e-010 ua=-9.840109e-010             lua=3.4853384e-016             wua=3.6060526e-017 pua=-1.1365577e-022            ub=1.8396323e-018             lub=1.5416072e-025 wub=1.7672762e-026             pub=-8.4171752e-032            uc=5.2213345e-010 luc=-3.7303514e-016            wuc=-1.902972e-017             puc=2.0562336e-023 vsat=99777.778                  wvsat=0.0055813333               a0=0.4510403 la0=3.7638193e-007             wa0=2.0972911e-007             pa0=-2.0550236e-013 ags=1.8611222                  lags=1.1543622e-006             wags=-2.396484e-007 pags=1.5627691e-013             keta=-0.03139326                lketa=-1.1817848e-007 wketa=2.8173719e-008             pketa=-1.8742515e-014            pclm=0.50222222 wpclm=-5.5813333e-008            pdiblc2=0.0010282066               lpdiblc2=-2.5374678e-010 wpdiblc2=-2.144052e-011             ppdiblc2=1.9287892e-016             aigbacc=0.010732107 laigbacc=-1.4556631e-009            waigbacc=1.6309114e-011             paigbacc=3.441863e-017 aigc=0.0096201292               laigc=2.326935e-011              waigc=6.723114e-011 paigc=-1.7228449e-017            bigc=0.00093700444              wbigc=5.5143573e-011 aigsd=0.0095473107               laigsd=-1.3123459e-010            waigsd=-2.3288372e-011 paigsd=5.530808e-017              bigsd=0.00058                    tvoff=0.0022527 ltvoff=-5.13073e-010              wtvoff=-1.22165e-010              ptvoff=1.34471e-016 kt1=-0.1056463                 lkt1=2.6995428e-012             wkt1=-2.611934e-009 pkt1=-1.1696846e-018            kt2=-0.031687771               lkt2=-2.5815003e-013 wkt2=-2.8933608e-009            pkt2=-2.204961e-020             ute=-0.675 ua1=2.7096952e-009             lua1=1.1397495e-016             wua1=7.1097192e-017 pua1=-6.2229291e-023            ub1=-2.3040136e-018            lub1=-1.7801467e-030 wub1=-6.7969585e-026            pub1=9.7196012e-037             uc1=-3.7103706e-010 luc1=9.1550215e-017             wuc1=1.3551396e-016             puc1=-4.9986468e-023 at=150000                     wat=0                          lcit=-8.3956196e-011 wcit=-4.8257867e-010            pcit=4.5840083e-017             lu0=2.1082351e-009 pu0=-1.1510964e-015            lvsat=0                          pvsat=0 lpclm=0                          ppclm=0                          lat=0 pat=0                          leta0=0                          peta0=0 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00166856                 lvoff_mcl=2.98496e-09                wvoff_mcl=2.67e-15 pvoff_mcl=-2.1e-21 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.16 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.59068068 lvth0=-3.3440538e-010            wvth0=-3.1006254e-009            pvth0=1.4849392e-015 k2=-0.049577176               lk2=-3.9219411e-009            wk2=7.4394616e-010 pk2=3.9030399e-016             cit=0.0067296256               voff=-0.20570651 lvoff=-5.1738129e-009            wvoff=1.884974e-009              pvoff=4.1511079e-016 eta0=0.022963911                weta0=1.9612805e-009             etab=-0.0128608 wetab=-3.8980032e-009            u0=0.043360072                wu0=-3.2111455e-009 ua=-1.4570843e-010            lua=-4.0258518e-016            wua=-1.6015114e-016 pua=6.2149883e-023             ub=2.2394903e-018             lub=-2.0411202e-025 wub=-1.2597145e-025            pub=4.4533461e-032             uc=1.3136983e-010 luc=-2.2910946e-017            wuc=7.8037927e-018             puc=-3.4804915e-024 vsat=94367.633                  wvsat=0.0085352726               a0=0.68371916 la0=1.6790167e-007             wa0=1.822761e-007              pa0=-1.8090446e-013 ags=2.8967678                  lags=2.2642379e-007             wags=-1.9250143e-008 pags=-4.119993e-014             keta=-0.21318737                lketa=4.4709038e-008 wketa=2.7319287e-008             pketa=-1.7976944e-014            pclm=0.58416861 wpclm=-1.5467073e-007            pdiblc2=0.00089031101              lpdiblc2=-1.3019231e-010 wpdiblc2=-5.2182986e-011            ppdiblc2=2.2042417e-016             aigbacc=0.0095569272 laigbacc=-4.0270157e-010            waigbacc=4.5606597e-011             paigbacc=8.1680851e-018 aigc=0.0091804541               laigc=4.1721823e-010             waigc=1.8778241e-010 paigc=-1.2524239e-016            bigc=0.00037535279              wbigc=2.1915911e-010 aigsd=0.0094273258               laigsd=-2.3728119e-011            waigsd=3.3562044e-011 paigsd=4.3701074e-018             bigsd=0.00068462169              wbigsd=-2.8875586e-011 tvoff=0.00182202                 ltvoff=-1.2718e-010               wtvoff=7.00051e-012 ptvoff=1.87383e-017               kt1=-0.10295556                lkt1=-2.408203e-009 wkt1=-2.6899517e-009            pkt1=6.873418e-017              kt2=-0.0140344 lkt2=-1.5817679e-008            wkt2=-2.6756757e-009            pkt2=-1.9506784e-016 ute=-0.64819485                wute=-3.872205e-010             ua1=3.3514238e-009 lua1=-4.610139e-016             wua1=8.1395205e-017             pua1=-7.1456311e-023 ub1=-2.2313351e-018            lub1=-6.5121668e-026            wub1=-3.341219e-025 pub1=2.3847344e-031             uc1=-5.2943459e-010            luc1=2.334744e-016 wuc1=9.1463681e-017             puc1=-1.0517417e-023            at=84624.109 wat=0.054972546                lcit=-1.7109864e-009            wcit=-1.0249525e-009 pcit=5.3180708e-016             lu0=-7.2324079e-009            pu0=1.3771579e-015 lvsat=0.0048474901               pvsat=-2.6467296e-009            lpclm=-7.3423964e-008 ppclm=8.8576226e-014             lbigc=5.0323988e-010             pbigc=-1.4695793e-016 lbigsd=-9.3741033e-011            pbigsd=2.5872525e-017             lute=-2.4017415e-008 pute=3.4694957e-016             lat=0.058576798                pat=-4.9255401e-008 leta0=0                          peta0=0                          jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499999 lvoff_mcl=-8.4e-15                   wvoff_mcl=-7e-16                     pvoff_mcl=1.2e-21 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.17 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.59210678 lvth0=-9.7044904e-010            wvth0=2.0693433e-009             pvth0=-8.2086687e-016 k2=-0.046063741               lk2=-5.4889329e-009            wk2=-1.4218914e-010 pk2=7.8552033e-016             cit=0.0014236277               voff=-0.21326431 lvoff=-1.8030353e-009            wvoff=4.9318188e-009             pvoff=-9.4378198e-016 eta0=0.018268504                weta0=4.524973e-009              etab=-0.0128608 wetab=-3.8980032e-009            u0=0.032113529                wu0=-4.2674302e-010 ua=-9.2225457e-010            lua=-5.62456e-017              wua=-9.8298347e-018 pua=-4.8934204e-024            ub=2.157682e-018              lub=-1.6762552e-025 wub=-7.2641292e-026            pub=2.0748211e-032             uc=2.1850546e-010 luc=-6.1773436e-017            wuc=-1.3347342e-017            puc=5.9529147e-024 vsat=94668.606                  wvsat=0.0054029413               a0=2.1843665 la0=-5.0138702e-007            wa0=-4.4085064e-007            pa0=9.7010063e-014 ags=3.3078063                  lags=4.3100627e-008             wags=4.0071111e-008 pags=-6.7657209e-014            keta=-0.17673274                lketa=2.8450275e-008 wketa=8.6190575e-009             pketa=-9.6366418e-015            pclm=0.2020917 wpclm=7.361793e-008              pdiblc2=-0.00067142564             lpdiblc2=5.6634224e-010 wpdiblc2=8.4252373e-010             ppdiblc2=-1.7861503e-016            aigbacc=0.0090875353 laigbacc=-1.9335276e-010            waigbacc=7.4073558e-011             paigbacc=-4.5281797e-018 aigc=0.0097634837               laigc=1.5718702e-010             waigc=-4.5667152e-011 paigc=-2.1123882e-017            bigc=0.0010528803               wbigc=-3.5353692e-011 aigsd=0.0093210194               laigsd=2.3684527e-011             waigsd=7.1297199e-011 paigsd=-1.2459772e-017            bigsd=0.00034657561              wbigsd=7.3126916e-011 tvoff=0.00219859                 ltvoff=-2.95132e-010              wtvoff=-1.10006e-010 ptvoff=7.0923e-017                kt1=-0.067663833               lkt1=-1.8148313e-008 wkt1=-1.8218493e-008            pkt1=6.9944638e-015             kt2=-0.056781693 lkt2=3.2476137e-009             wkt2=-6.9067522e-009            pkt2=1.6919923e-015 ute=-0.28534234                wute=-1.2102821e-007            ua1=2.0391848e-009 lua1=1.242447e-016              wua1=2.9886634e-016             pua1=-1.6844844e-022 ub1=-1.2652199e-018            lub1=-4.9600908e-025            wub1=-3.7306209e-025 pub1=2.5584077e-031             uc1=3.1330713e-010             luc1=-1.423884e-016 wuc1=1.9775436e-017             puc1=2.145554e-023              at=284878.92 wat=-0.088455338               lcit=6.554887e-010              wcit=6.7309926e-010 pcit=-2.2552403e-016            lu0=-2.2164497e-009            pu0=1.3531442e-016 lvsat=0.0047132561               pvsat=-1.2497098e-009            lpclm=9.6982337e-008 ppclm=-1.3240516e-014            lbigc=2.0106263e-010             pbigc=-3.3445214e-017 lbigsd=5.7027517e-011             pbigsd=-1.9620591e-017            lute=-1.8584963e-007 pute=5.415283e-014              lat=-0.030736846               pat=1.4713435e-008 leta0=2.0941517e-009             peta0=-1.1434068e-015 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00499999                 lvoff_mcl=1.6e-15                    wvoff_mcl=3.7e-15 pvoff_mcl=1e-22                      u0_ff=-0.00054963                u0_fs=-0.00036642 wu0_ff=1.51698e-10                wu0_fs=1.01132e-10                lu0_ff=2.45135e-10 lu0_fs=1.63423e-10                pu0_ff=-6.76572e-17               pu0_fs=-4.51048e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.18 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.60730559 lvth0=-4.1925957e-009            wvth0=-3.6606412e-009            pvth0=3.9388985e-016 k2=-0.069204846               lk2=-5.8301856e-010            wk2=2.7928048e-009 pk2=1.6330162e-016             cit=0.0050534253               voff=-0.2113606 lvoff=-2.2066223e-009            wvoff=-1.6181125e-009            pvoff=4.4480344e-016 eta0=0.033085071                weta0=-2.9850034e-009            etab=-0.0128608 wetab=-3.8980032e-009            u0=0.02365126                 wu0=-1.2293994e-010 ua=-1.0954754e-009            lua=-1.9522776e-017            wua=-7.4223022e-017 pua=8.7579352e-024             ub=1.4817729e-018             lub=-2.4332807e-026 wub=4.9874972e-026             pub=-5.2252372e-033            uc=-3.6075583e-011 luc=-7.8022545e-018            wuc=7.5150181e-018             puc=1.5300943e-024 vsat=130421.87                  wvsat=-0.0048930088              a0=2.9873792 la0=-6.7162572e-007            wa0=-3.527757e-007             pa0=7.8338177e-014 ags=3.5111111                  lags=0                          wags=-2.7906667e-007 pags=0                          keta=0.05201358                 lketa=-2.0043946e-008 wketa=-6.2931748e-008            pketa=5.532129e-015              pclm=0.44648183 wpclm=2.4838705e-008             pdiblc2=0.002                      aigbacc=0.0086487176 laigbacc=-1.0032341e-010            waigbacc=4.661671e-011              paigbacc=1.292672e-018 aigc=0.010636011                laigc=-2.7788688e-011            waigc=-1.5555255e-010 paigc=2.1718218e-018             bigc=0.0021822059               wbigc=-2.1821862e-010 aigsd=0.0094995581               laigsd=-1.4165669e-011            waigsd=2.2028977e-011 paigsd=-2.0149088e-018            bigsd=0.00056727682              wbigsd=4.6245333e-013 tvoff=0.00074024                 ltvoff=1.40387e-011               wtvoff=1.47599e-010 ptvoff=1.63109e-017               kt1=-0.20180214                lkt1=1.0289008e-008 wkt1=1.6991906e-008             pkt1=-4.7014082e-016            kt2=-0.050660505 lkt2=1.9499219e-009             wkt2=4.2555566e-009             pkt2=-6.7441717e-016 ute=-1.4563174                 wute=2.1877826e-007             ua1=4.3520396e-009 lua1=-3.6608053e-016            wua1=-6.2131704e-016            pua1=2.6630439e-023 ub1=-6.0767656e-018            lub1=5.2403861e-025             wub1=1.1114795e-024 pub1=-5.8882043e-032            uc1=-7.1090796e-010            luc1=7.4745196e-017 wuc1=1.7307917e-016             puc1=-1.1044851e-023            at=211361.29 wat=-0.032073124               lcit=-1.1402838e-010            wcit=-7.5890353e-010 pcit=7.8060561e-017             lu0=-4.2244862e-010            pu0=7.0908165e-017 lvsat=-0.0028664364              pvsat=9.330316e-010              lpclm=4.5171629e-008 ppclm=-2.8993202e-015            lbigc=-3.8354404e-011            pbigc=5.3221504e-018 lbigsd=1.023886e-011              pbigsd=-4.2157246e-018            lute=6.2397075e-008 pute=-1.788614e-014             lat=-0.015151109               pat=2.7604057e-009 leta0=-1.0469605e-009            peta0=4.4870816e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00499999                 lvoff_mcl=1.34e-15                   wvoff_mcl=-7e-16 pvoff_mcl=4e-23                      u0_ff=0.000606666                u0_fs=0.000680494 wu0_ff=-1.6744e-10                wu0_fs=-1.87816e-10               ua1_ff=1.39541e-11 lua1_ff=-2.95828e-18               wua1_ff=-7.61896e-18               pua1_ff=1.61522e-24 lu0_ff=4e-18                      lu0_fs=-5.85225e-11               pu0_ff=-2e-24 pu0_fs=1.61522e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.19 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.56510829 lvth0=-5.6362793e-010            wvth0=-7.0396995e-009            pvth0=6.8448886e-016 k2=-0.081923521               lk2=5.1078746e-010             wk2=7.273364e-009 pk2=-2.2202647e-016            cit=0.0022741782               voff=-0.24796361 lvoff=9.4123702e-010             wvoff=1.2144143e-008             pvoff=-7.3875053e-016 eta0=0.0096765432               weta0=5.3332741e-009             etab=-0.0041010778 wetab=-1.0316536e-008            u0=0.016915517                wu0=1.2581566e-009 ua=-2.169523e-009             lua=7.2845316e-017             wua=1.7095403e-016 pua=-1.2327291e-023            ub=1.9573222e-018             lub=-6.5230044e-026 wub=-1.4246353e-025            pub=1.1315874e-032             uc=-1.1818073e-010 luc=-7.412115e-019             wuc=5.5546592e-017             puc=-2.6006211e-024 vsat=75335.19                   wvsat=0.0057016529               a0=-1.2664089 la0=-3.0579995e-007            wa0=1.2950926e-006             pa0=-6.3378496e-014 ags=3.5111111                  lags=0                          wags=-2.7906667e-007 pags=0                          keta=-0.080145062               lketa=-8.6783025e-009 wketa=1.3410704e-008             pketa=-1.0333218e-015            pclm=1.3621037 wpclm=2.0557911e-009             pdiblc2=0.002                      aigbacc=0.0068545353 laigbacc=5.3976263e-011             waigbacc=1.440549e-010              paigbacc=-7.0870126e-018 aigc=0.010683972                laigc=-3.1913351e-011            waigc=-3.8475615e-010 paigc=2.1883332e-017             bigc=0.0020464374               wbigc=-4.7563192e-010 aigsd=0.0095316358               laigsd=-1.6924357e-011            waigsd=-1.248893e-010 paigsd=1.0620063e-017             bigsd=0.0011616111               wbigsd=-2.5088093e-010 tvoff=-0.000849068               ltvoff=1.50719e-010               wtvoff=7.90942e-010 ptvoff=-3.90166e-017              kt1=-0.12343609                lkt1=3.5495273e-009 wkt1=1.0273962e-008             pkt1=1.076023e-016              kt2=-0.023055552 lkt2=-4.2410407e-010            wkt2=-5.5371351e-009            pkt2=1.6775432e-016 ute=-0.80822833                wute=2.5799713e-008             ua1=4.5961031e-010 lua1=-3.1331608e-017            wua1=-4.6501873e-017            pua1=-2.2803665e-023 ub1=-3.503921e-019             lub1=3.1570494e-026             wub1=1.0277715e-025 pub1=2.7866357e-032             uc1=-9.8366599e-011            luc1=2.2066639e-017 wuc1=5.4135848e-017             puc1=-8.157256e-025             at=24729.824 wat=0.0049477288               lcit=1.2498687e-010             wcit=2.6874701e-010 pcit=-1.0317385e-017            lu0=1.5682525e-010             pu0=-4.7866135e-017 lvsat=0.0018710183               pvsat=2.189069e-011              lpclm=-3.3571852e-008 ppclm=-9.3998956e-016            lbigc=-2.6678315e-011            pbigc=2.7459695e-017 lbigsd=-4.0873889e-011            pbigsd=1.7399807e-017             lute=6.6614167e-009 pute=-1.2899857e-015            lat=0.00089919689              pat=-4.2338764e-010 leta0=9.6617284e-010             peta0=-2.666637e-016             letab=-7.5333611e-010 petab=5.5199387e-016             jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499999 lvoff_mcl=-3.83e-15                  wvoff_mcl=4.1e-15                    pvoff_mcl=6.3e-22 u0_ff=0.00144926                 wu0_ff=-3.99996e-10               ua1_ff=-4.88395e-11 lua1_ff=2.44198e-18                wua1_ff=2.66664e-17                pua1_ff=-1.33332e-24 lu0_ff=-7.2463e-11                pu0_ff=1.99998e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.20 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.47326535 lvth0=4.0285191e-009             wvth0=2.9322472e-008             pvth0=-1.1336197e-015 k2=-0.10851874                lk2=1.8405485e-009             wk2=1.7806558e-008 pk2=-7.4868615e-016            cit=0.0036530554               voff=-0.11512133 lvoff=-5.700877e-009             wvoff=-3.3004169e-008            pvoff=1.5186651e-015 eta0=0.030649356                weta0=-9.2565555e-009            etab=-0.029530272 wetab=5.0928116e-009             u0=0.0079467481               wu0=5.9104055e-009 ua=-1.4667143e-009            lua=3.770488e-017              wua=-1.0997335e-016 pua=1.719078e-024              ub=7.2435522e-019             lub=-3.5816942e-027 wub=4.1354623e-025             pub=-1.6484614e-032            uc=-6.1729924e-010 luc=2.4214714e-017             wuc=1.0247127e-016             puc=-4.9468552e-024 vsat=-52230.275                 wvsat=0.053041623                a0=-17.14246 la0=4.8800261e-007             wa0=6.7665307e-006             pa0=-3.369504e-013 ags=3.5111111                  lags=0                          wags=-2.7906667e-007 pags=0                          keta=-0.63012895                lketa=1.8820892e-008 wketa=6.3131585e-008             pketa=-3.5193659e-015            pclm=1.2540107 wpclm=5.4093042e-008             pdiblc2=0.002                      aigbacc=0.0081995622 laigbacc=-1.3275081e-011            waigbacc=1.3464587e-010             paigbacc=-6.6165611e-018 aigc=0.010100852                laigc=-2.7573376e-012            waigc=4.2609584e-010 paigc=-1.8659268e-017            bigc=0.0012647034               wbigc=5.7709359e-010 aigsd=0.0086732964               laigsd=2.5992614e-011             waigsd=2.0391487e-010 paigsd=-5.8201453e-018            bigsd=-0.00028807767             wbigsd=3.1536064e-010 tvoff=-0.000349503               ltvoff=1.25741e-010               wtvoff=6.70947e-010 ptvoff=-3.30169e-017              kt1=-0.45777776                lkt1=2.0266611e-008 wkt1=1.0283781e-007             pkt1=-4.52059e-015              kt2=0.014959115 lkt2=-2.3248374e-009            wkt2=-1.8424333e-008            pkt2=8.1211423e-016 ute=-0.675                     ua1=1.4063132e-008             lua1=-7.1150769e-016 wua1=-3.755404e-015             pua1=1.6264144e-022             ub1=-1.7429808e-017 lub1=8.8554128e-025             wub1=4.7610758e-024             pub1=-2.0504857e-031 uc1=-1.6460185e-009            luc1=9.9449231e-017             wuc1=6.1973894e-016 puc1=-2.909588e-023             at=206208.9                   wat=-0.04126302 lcit=5.6043007e-011             wcit=1.25189e-009               pcit=-5.9474537e-017 lu0=6.052637e-010              pu0=-2.8047858e-016            lvsat=0.0082492915 pvsat=-2.3451078e-009            lpclm=-2.8167203e-008            ppclm=-3.5418521e-015 lbigc=1.2408384e-011             pbigc=-2.5176581e-017            lbigsd=3.161055e-011 pbigsd=-1.0912272e-017            lat=-0.0081747567              pat=1.8871498e-009 leta0=-8.2467785e-011            peta0=4.6282778e-016             letab=5.1812358e-010 petab=-2.1847354e-016            jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               voff_mcl=0.00499995 lvoff_mcl=-7.5e-15                   wvoff_mcl=-3.7e-14                   pvoff_mcl=-1.5e-22 ua1_fs=-9.11112e-11               lua1_fs=4.55556e-18                wua1_fs=-4.8e-23 pua1_fs=-2.6e-30 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.21 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.50142867 lvth0=2.8738231e-009             wvth0=-1.6866866e-009            pvth0=1.3775578e-016 k2=-0.028482622               lk2=-1.4409324e-009            wk2=-1.1605093e-008 pk2=4.5719151e-016             cit=0.00049240138              voff=-0.22399643 lvoff=-1.2369979e-009            wvoff=1.3278813e-008             pvoff=-3.7893719e-016 eta0=-0.01895059                weta0=1.124103e-008              etab=-0.028403334 wetab=-4.2655334e-009            u0=0.01611218                 wu0=-5.1424842e-010 ua=-8.1086485e-010            lua=1.0815053e-017             wua=-4.2027156e-016 pua=1.4441305e-023             ub=7.2059105e-019             lub=-3.4273632e-027 wub=3.8894781e-025             pub=-1.5476078e-032            uc=-9.5060385e-011 luc=2.8029208e-018             wuc=1.815289e-017              puc=-1.4898015e-024 vsat=88154.739                  wvsat=-0.014932775               a0=4.6005578 la0=-4.0346112e-007            wa0=-3.8454841e-006            pa0=9.8142205e-014 ags=3.5111111                  lags=0                          wags=-2.7906667e-007 pags=0                          keta=0.16502574                 lketa=-1.378045e-008 wketa=-6.4004328e-009            pketa=-6.6855319e-016            pclm=1.4892632 wpclm=-1.7114725e-007            pdiblc2=0.002                      aigbacc=0.0075638216 laigbacc=1.2790283e-011             waigbacc=-8.0180454e-011            paigbacc=2.1913183e-018 aigc=0.013355329                laigc=-1.3619092e-010            waigc=-5.8263104e-010 paigc=2.2698534e-017             bigc=0.0055449558               wbigc=-8.9671794e-010 aigsd=0.0083925905               laigsd=3.7501557e-011             waigsd=2.5006015e-010 paigsd=-7.7121017e-018            bigsd=-0.00027473715             wbigsd=2.2416825e-010 tvoff=0.0026344                  ltvoff=3.40083e-012               wtvoff=2.18912e-012 ptvoff=-5.5978e-018               kt1=-0.00024126838             lkt1=1.5076149e-009 wkt1=-1.0783674e-008            pkt1=1.3789077e-016             kt2=-0.079184293 lkt2=1.5350423e-009             wkt2=4.4787922e-010             pkt2=3.8353512e-017 ute=-0.57467091                wute=1.9310917e-007             ua1=-3.3541763e-009 lua1=2.6019503e-018             wua1=1.1709045e-015             pua1=-3.9337209e-023 ub1=5.2996163e-018             lub1=-4.6365108e-026            wub1=-1.3700685e-024 pub1=4.6328341e-032             uc1=2.1122805e-009             luc1=-5.4641027e-017 wuc1=-3.7979922e-016            puc1=1.1885184e-023             at=-26514.307 wat=0.012391165                lcit=1.8562982e-010             wcit=-1.5005694e-009 pcit=5.3376302e-017             lu0=2.7048099e-010             pu0=-1.7067771e-017 lvsat=0.0024935059               pvsat=4.4184252e-010             lpclm=-3.7812553e-008 ppclm=5.6929997e-015             lbigc=-1.6308196e-010            pbigc=3.5249692e-017 lbigsd=3.1063589e-011             pbigsd=-7.1733841e-018            lute=-4.1134925e-009 pute=-7.9174761e-015            lat=0.0013668946               pat=-3.1267176e-010 leta0=1.95113e-009               peta0=-3.7757321e-016            letab=4.7191916e-010 petab=1.6521861e-016             jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               vth0_mc=-0.0181728 lvth0_mc=7.45086e-10                wvth0_mc=9.92237e-09                pvth0_mc=-4.06817e-16 voff_ff=-0.00711106                voff_ss=0.0143802                  voff_mcl=0.00499994 voff_mc=-0.0181728                 lvoff_ff=2.91555e-10                lvoff_ss=-5.8959e-10 lvoff_mcl=-4.42e-15                  lvoff_mc=7.45086e-10                wvoff_ff=1.9e-15 wvoff_ss=-3.96895e-09               wvoff_mcl=3.96e-14                   wvoff_mc=9.92237e-09 pvoff_ff=-1.3e-22                   pvoff_ss=1.62727e-16                pvoff_mcl=1.9e-22 pvoff_mc=-4.06817e-16               u0_mc=-0.00173827                wu0_mc=-9.92241e-10 ua_ff=7.90158e-13                lua_ff=-3.23957e-20               wua_ff=-1.98448e-17 pua_ff=8.13635e-25                vsat_ff=10785.2                    vsat_fs=-3555.55 vsat_mc=-7585.18                   wvsat_ff=-0.00297671                wvsat_fs=-4.1e-09 wvsat_mc=0.0119068                  ua1_fs=9.11112e-11                lua1_fs=-2.91555e-18 wua1_fs=4.8e-23                    pua1_fs=1.3e-30                    lu0_mc=7.12691e-11 pu0_mc=4.06818e-17                lvsat_ff=-0.000442193               lvsat_fs=0.000145778 lvsat_mc=0.000310993                pvsat_ff=1.22045e-10                pvsat_fs=3.7e-17 pvsat_mc=-4.8818e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.22 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.54914254 lvth0=1.5418521e-008             wvth0=5.7009416e-009             pvth0=-4.7685783e-016 k2=-0.049030028               lk2=-9.4265562e-009            wk2=3.2119009e-010 pk2=2.1530598e-015             cit=0.0035734571               voff=-0.20396435 lvoff=-1.3974636e-008            wvoff=2.8003315e-009             pvoff=1.5931482e-015 eta0=0.040674815                weta0=-2.9269289e-009            etab=-0.028380148 wetab=3.8533689e-010             u0=0.031483611                wu0=1.1218637e-011 ua=-8.8177146e-010            lua=-5.6091798e-018            wua=7.84244e-018 pua=-1.5912299e-023            ub=1.8995054e-018             lub=-2.3557701e-025 wub=1.1477928e-027             pub=2.3395862e-032             uc=5.3368124e-010 luc=-3.7696358e-016            wuc=-2.2216912e-017            puc=2.1646584e-023 vsat=112962.96                  wvsat=0.0019422222               a0=0.80708022 la0=-1.7334159e-007            wa0=1.114621e-007              pa0=-5.377867e-014 ags=0.82745016                 lags=2.1670777e-006             wags=4.5645086e-008 pags=-1.2323256e-013            keta=0.051762746                lketa=-1.7209486e-007 wketa=5.2226615e-009             pketa=-3.861596e-015             pclm=0.3 wpclm=0                          pdiblc2=0.0010161623               lpdiblc2=-1.4539567e-010 wpdiblc2=-1.8116275e-011            ppdiblc2=1.6297401e-016             aigbacc=0.010588578 laigbacc=-1.3694864e-009            waigbacc=5.5923153e-011             paigbacc=1.0633856e-017 aigc=0.010069877                laigc=-4.0319087e-011            waigc=-5.6899144e-011 paigc=3.2196009e-019             bigc=0.0012990178               wbigc=-4.4772107e-011 aigsd=0.0094022829               laigsd=1.3305017e-010             waigsd=1.6739287e-011 paigsd=-1.7634514e-017            bigsd=0.00062036727              wbigsd=-1.1141368e-011 tvoff=0.00161923                 ltvoff=-2.91792e-010              wtvoff=5.26744e-011 ptvoff=7.33971e-017               kt1=-0.11662991                lkt1=-8.3047716e-013 wkt1=4.1954172e-010             pkt1=-1.9539908e-019            kt2=-0.046344634 lkt2=-2.922426e-013             wkt2=1.1519334e-009             pkt2=-1.2640059e-020 ute=-0.63822463                wute=-1.0150002e-008            ua1=3.6106421e-009 lua1=-1.8133152e-016            wua1=-1.7756416e-016            pua1=1.9275296e-023 ub1=-3.3737613e-018            lub1=1.4403341e-030             wub1=2.2728078e-025 pub1=8.3107422e-038             uc1=7.3316872e-012             luc1=-1.5258401e-016 wuc1=3.1084188e-017             puc1=1.7394577e-023             at=150000 wat=0                          lcit=-3.1450746e-010            wcit=-1.1265957e-010 pcit=1.0947223e-016             lu0=-3.6022274e-009            pu0=4.249913e-016 lvsat=0                          pvsat=0                          lpclm=0 ppclm=0                          lbigsd=-1.3094951e-016            pbigsd=3.6142065e-023 lute=1.6841368e-012             pute=-4.6482175e-019            lat=0 pat=0                          leta0=0                          peta0=0 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' vth0_mc=0.000388729                lvth0_mc=-3.50089e-09               wvth0_mc=-1.07289e-10 pvth0_mc=9.66247e-16                voff_ff=0.000233237                voff_mcl=0.00166856 voff_mc=0.000777458                lvoff_ff=-2.10054e-09               lvoff_mcl=2.98498e-09 lvoff_mc=-7.00179e-09               wvoff_ff=-6.43735e-11               wvoff_mcl=-2.2e-16 wvoff_mc=-2.14578e-10               pvoff_ff=5.79748e-16                pvoff_mcl=-3.1e-22 pvoff_mc=1.93249e-15                ags_ff=-0.0194365                 ags_ss=0.0116619 lags_ff=1.75045e-07                lags_ss=-1.05027e-07               wags_ff=5.36446e-09 wags_ss=-3.21868e-09               pags_ff=-4.83123e-14               pags_ss=2.89874e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.23 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.5518118 lvth0=1.3026862e-008             wvth0=7.6271834e-009             pvth0=-2.2027705e-015 k2=-0.057578296               lk2=-1.767308e-009             wk2=2.9522555e-009 pk2=-2.0437474e-016            cit=0.0025986315               voff=-0.21684749 lvoff=-2.4313395e-009            wvoff=4.9598852e-009             pvoff=-3.4181186e-016 eta0=0.040674815                weta0=-2.9269289e-009            etab=-0.028380148 wetab=3.8533689e-010             u0=0.028222724                wu0=9.6676266e-010 ua=-7.3715394e-010            lua=-1.3518647e-016            wua=3.0878191e-018 pua=-1.1652159e-023            ub=1.5855124e-018             lub=4.5760658e-026 wub=5.4526433e-026             pub=-2.4431399e-032            uc=1.7520474e-010 luc=-5.5768633e-017            wuc=-4.2946418e-018            puc=5.5882301e-024 vsat=121979.87                  wvsat=0.00091429464              a0=1.069738 la0=-4.0868293e-007            wa0=7.5734911e-008             pa0=-2.1767112e-014 ags=3.1412158                  lags=9.3943664e-008             wags=-8.6717805e-008 pags=-4.6354145e-015            keta=-0.068625939               lketa=-6.4226596e-008 wketa=-1.2579668e-008            pketa=1.2089291e-014             pclm=0.010446155 wpclm=3.6766698e-009             pdiblc2=-0.00076383655             lpdiblc2=1.4494833e-009 wpdiblc2=4.0436174e-010             ppdiblc2=-2.1556629e-016            aigbacc=0.0094328184 laigbacc=-3.3392543e-010            waigbacc=7.9860636e-011             paigbacc=-1.0814129e-017 aigc=0.010067128                laigc=-3.7856397e-011            waigc=-5.6939602e-011 paigc=3.5821073e-019             bigc=0.0012884114               wbigc=-3.2845067e-011 aigsd=0.0095324829               laigsd=1.6391014e-011             waigsd=4.5386839e-012 paigsd=-6.7027733e-018            bigsd=0.0005794714               wbigsd=1.4589263e-013 tvoff=0.00122083                 ltvoff=6.51744e-011               wtvoff=1.7293e-010 ptvoff=-3.43515e-017              kt1=-0.11354398                lkt1=-2.7658206e-009 wkt1=2.3245237e-010             pkt1=1.6743666e-016             kt2=-0.023127806 lkt2=-2.080257e-008             wkt2=-1.6589555e-010            pkt2=1.1807621e-015 ute=-0.78357523                wute=3.6977764e-008             ua1=3.9899085e-009 lua1=-5.2115419e-016            wua1=-9.4826566e-017            pua1=-5.4857591e-023 ub1=-4.5227145e-018            lub1=1.0294636e-024             wub1=2.9829882e-025 pub1=-6.3632081e-032            uc1=-5.6234403e-010            luc1=3.5784544e-016 wuc1=1.0054669e-016             puc1=-4.4843822e-023            at=325697.88 wat=-0.011563814               lcit=5.5893627e-010             wcit=1.1520181e-010 pcit=-9.4691563e-017            lu0=-6.804728e-010             pu0=-4.3117614e-016 lvsat=-0.0080791501              pvsat=9.2102312e-010             lpclm=2.5944025e-007 ppclm=-3.2942962e-015            lbigc=9.5032961e-012             pbigc=-1.0686628e-017 lbigsd=3.6642569e-011             pbigsd=-1.0113349e-017            lute=1.3023582e-007 pute=-4.2226943e-014            lat=-0.1574253                 pat=1.0361178e-008 leta0=0                          peta0=0                          jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)' jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               vth0_mc=-0.00700576 lvth0_mc=3.12457e-09                wvth0_mc=1.93359e-09                pvth0_mc=-8.62381e-16 voff_ff=-0.00420346                voff_mcl=0.00499998                 voff_mc=-0.0140115 lvoff_ff=1.87474e-09                lvoff_mcl=5e-16                      lvoff_mc=6.24914e-09 wvoff_ff=1.16015e-09                wvoff_mcl=-1e-17                     wvoff_mc=3.86718e-09 pvoff_ff=-5.17429e-16               pvoff_mcl=2e-22                      pvoff_mc=-1.72476e-15 ags_ff=0.350288                   ags_ss=-0.210173                  lags_ff=-1.56228e-07 lags_ss=9.37371e-08                wags_ff=-9.66795e-08               wags_ss=5.80077e-08 pags_ff=4.31191e-14                pags_ss=-2.58714e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.24 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.59080042 lvth0=-4.3620618e-009            wvth0=2.4298993e-009             pvth0=1.1521824e-016 k2=-0.053263445               lk2=-3.6917315e-009            wk2=1.8449293e-009 pk2=2.8949272e-016             cit=0.0054255777               voff=-0.19873421 lvoff=-1.0509863e-008            wvoff=9.2151222e-010             pvoff=1.4593025e-015 eta0=0.048500494                weta0=-3.8190563e-009            etab=-0.028380148 wetab=3.8533689e-010             u0=0.031801409                wu0=-3.405977e-010 ua=-8.3827854e-010            lua=-9.0084902e-017            wua=-3.3007217e-017 pua=4.4462271e-024             ub=1.9024167e-018             lub=-9.5578633e-026 wub=-2.188071e-027             pub=8.6326964e-034             uc=1.7683734e-010 luc=-5.6496773e-017            wuc=-1.8469413e-018            puc=4.4965557e-024 vsat=104432.35                  wvsat=0.0027081481               a0=0.54137156 la0=-1.7303151e-007            wa0=1.2615955e-008             pa0=6.383942e-015 ags=3.8048433                  lags=-2.0203419e-007            wags=-9.7111111e-008 pags=1.7504824e-028             keta=-0.21011707                lketa=-1.1215516e-009 wketa=1.7833132e-008             pketa=-1.4748177e-015            pclm=0.5390692 wpclm=-1.938786e-008             pdiblc2=0.0026077759               lpdiblc2=-5.4255907e-011 wpdiblc2=-6.2535904e-011            ppdiblc2=-7.329944e-018             aigbacc=0.0091529628 laigbacc=-2.0910985e-010            waigbacc=5.6015558e-011             paigbacc=-1.7922419e-019 aigc=0.0098601087               laigc=5.4474264e-011             waigc=-7.2335629e-011 paigc=7.2248386e-018             bigc=0.0012015523               wbigc=-7.6387168e-011 aigsd=0.0097190285               laigsd=-6.680832e-011             waigsd=-3.8553305e-011 paigsd=1.2516254e-017             bigsd=0.00078833814              wbigsd=-4.8799543e-011 tvoff=0.00113079                 ltvoff=1.0533e-010                wtvoff=1.84708e-010 ptvoff=-3.96045e-017              kt1=-0.17083406                lkt1=2.2785554e-008 wkt1=1.0256489e-008             pkt1=-4.3032835e-015            kt2=-0.1000782 lkt2=1.3517305e-008             wkt2=5.0430833e-009             pkt2=-1.1424425e-015 ute=-0.5866286                 wute=-3.78732e-008              ua1=4.7549371e-009 lua1=-8.6235698e-016            wua1=-4.5068132e-016            pua1=1.0385363e-022 ub1=-4.1873398e-018            lub1=8.7988646e-025             wub1=4.3344303e-025 pub1=-1.239064e-031             uc1=3.1109577e-010             luc1=-3.1708714e-017 wuc1=2.0385772e-017             puc1=-9.0920543e-024            at=-89923.076 wat=0.014990012                lcit=-7.0188173e-010            wcit=-4.3143894e-010 pcit=1.4911021e-016             lu0=-2.2765662e-009            pu0=1.5190658e-016 lvsat=-0.00025295518             pvsat=1.2096448e-010             lpclm=2.3674366e-008 ppclm=6.9924841e-015             lbigc=4.8242472e-011             pbigc=8.7331496e-018 lbigsd=-5.6511997e-011            pbigsd=1.1716315e-017             lute=4.2397623e-008 pute=-8.8434126e-015            lat=0.027941647                pat=-1.4818288e-009 leta0=-3.4902528e-009            peta0=3.9788882e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00500005                 lvoff_mcl=7.9e-15                    wvoff_mcl=9.3e-16 pvoff_mcl=-7.1e-22 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.25 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.58570927 lvth0=-3.2827386e-009            wvth0=2.2999415e-009             pvth0=1.4276931e-016 k2=-0.07160794                lk2=1.9730133e-010             wk2=3.4560585e-009 pk2=-5.2066666e-017            cit=0.00061419128              voff=-0.25416031 lvoff=1.2404706e-009             wvoff=1.019461e-008              pvoff=-5.0659421e-016 eta0=0.027385656                weta0=-1.4119647e-009            etab=-0.028380148 wetab=3.8533689e-010             u0=0.020634481                wu0=7.0969106e-010 ua=-1.2833245e-009            lua=4.2648288e-018             wua=-2.2376695e-017 pua=2.1925563e-024             ub=1.5704904e-018             lub=-2.5210269e-026 wub=2.5388945e-026             pub=-4.9830577e-033            uc=-1.2013059e-010 luc=6.4604291e-018             wuc=3.0714201e-017             puc=-2.4064064e-024 vsat=97666.662                  wvsat=0.0041474291               a0=1.0721646 la0=-2.8555964e-007            wa0=1.7582352e-007             pa0=-2.8216062e-014 ags=2.8518519                  lags=0                          wags=-9.7111111e-008 pags=0                          keta=-0.26824104                lketa=1.1200729e-008 wketa=2.5458526e-008             pketa=-3.0914012e-015            pclm=0.45860127 wpclm=2.1493741e-008             pdiblc2=0.0023518519               wpdiblc2=-9.7111111e-011 aigbacc=0.0086350401               laigbacc=-9.9310227e-011            waigbacc=5.0391704e-011 paigbacc=1.0130328e-018             aigc=0.01033316                 laigc=-4.5812636e-011 waigc=-7.1965784e-011            paigc=7.1464315e-018             bigc=0.0016536035 wbigc=-7.2324348e-011            aigsd=0.0094958319               laigsd=-1.9490646e-011 waigsd=2.3057396e-011             paigsd=-5.4521497e-019            bigsd=0.00055182023 wbigsd=4.7284741e-012             tvoff=0.00146666                 ltvoff=3.41256e-011 wtvoff=-5.28933e-011              ptvoff=1.07669e-017               kt1=-0.085528814 lkt1=4.7008421e-009             wkt1=-1.5099533e-008            pkt1=1.072193e-015 kt2=-0.033820374               lkt2=-5.2935391e-010            wkt2=-3.9231961e-010 pkt2=9.8629553e-018             ute=-0.30702851                wute=-9.8425472e-008 ua1=1.7042057e-009             lua1=-2.1560192e-016            wua1=1.0948512e-016 pua1=-1.4901657e-023            ub1=-9.8992086e-019            lub1=2.0203363e-025 wub1=-2.9248967e-025            pub1=2.9991332e-032             uc1=4.3755706e-011 luc1=2.496738e-017              wuc1=-3.5208003e-017            puc1=2.6938261e-024 at=51150.95                   wat=0.012144931                lcit=3.1813219e-010 wcit=4.6632505e-010             pcit=-4.1215755e-017            lu0=9.0822413e-011 pu0=-7.0754642e-017            lvsat=0.0011813704               pvsat=-1.8416309e-010 lpclm=4.0733568e-008             ppclm=-1.6744153e-015            lbigc=-4.759238e-011 pbigc=7.8718316e-018             lbigsd=-6.3701989e-012            pbigsd=3.6837558e-019 lute=-1.6877596e-008            pute=3.9936688e-015             lat=-0.0019660466 pat=-8.786716e-010             leta0=9.8609289e-010             peta0=-1.1241459e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00499995                 lvoff_mcl=-4.04e-15                  wvoff_mcl=3.13e-15 pvoff_mcl=2.4e-22                    ua1_ff=-2.32569e-11               lua1_ff=4.93046e-18 wua1_ff=2.65129e-18                pua1_ff=-5.62073e-25 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.26 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.5274739 lvth0=1.7255032e-009             wvth0=3.3473906e-009             pvth0=5.2688688e-017 k2=-0.073604016               lk2=3.6896386e-010             wk2=4.9771805e-009 pk2=-1.8288315e-016            cit=0.0026267708               voff=-0.23432119 lvoff=-4.6569452e-010            wvoff=8.3788331e-009             pvoff=-3.5043742e-016 eta0=0.038851852                weta0=-2.7191111e-009            etab=-0.045953708 wetab=1.2347894e-009             u0=0.022689938                wu0=-3.3558363e-010 ua=-1.3586795e-009            lua=1.0745366e-017             wua=-5.2838775e-017 pua=4.8122952e-024             ub=1.3353298e-018             lub=-4.9864517e-027 wub=2.9206382e-026             pub=-5.3113574e-033            uc=5.7662911e-011 luc=-8.8298122e-018            wuc=7.0137461e-018             puc=-3.6816731e-025 vsat=84785.922                  wvsat=0.0030932508               a0=3.7493348 la0=-5.1579627e-007            wa0=-8.9252664e-008            pa0=-5.41951e-015 ags=2.8518519                  lags=0                          wags=-9.7111111e-008 pags=0                          keta=0.039674897                lketa=-1.5280041e-008 wketa=-1.9659605e-008            pketa=7.8875803e-016             pclm=1.5670561 wpclm=-5.4511056e-008            pdiblc2=0.0023518519               wpdiblc2=-9.7111111e-011 aigbacc=0.0069141122               laigbacc=4.8689571e-011             waigbacc=1.2761169e-010 paigbacc=-5.6278857e-018            aigc=0.0083275304               laigc=1.2667152e-010 waigc=2.656217e-010              paigc=-2.1886093e-017            bigc=-0.00076602212 wbigc=3.006069e-010              aigsd=0.0089134597               laigsd=3.0593359e-011 waigsd=4.5727296e-011             paigsd=-2.4948263e-018            bigsd=7.8252263e-005 wbigsd=4.8126109e-011             tvoff=0.00134848                 ltvoff=4.42893e-011 wtvoff=1.84419e-010               ptvoff=-9.64197e-018              kt1=-0.079539075 lkt1=4.1857245e-009             wkt1=-1.8416126e-009            pkt1=-6.7988106e-017 kt2=-0.030987933               lkt2=-7.7294381e-010            wkt2=-3.3477979e-009 pkt2=2.6403409e-016             ute=-0.26477911                wute=-1.2419227e-007 ua1=1.3453121e-009             lua1=-1.8473707e-016            wua1=-2.9095556e-016 pua1=1.9536242e-023             ub1=-1.0429611e-018            lub1=2.0659509e-025 wub1=2.939262e-025              pub1=-2.0440432e-032            uc1=1.4115226e-011 luc1=2.7516461e-017             wuc1=2.3090864e-017             puc1=-2.3198765e-024 at=33982.251                  wat=0.0023940592               lcit=1.4505035e-010 wcit=1.7143146e-010             pcit=-1.5854906e-017            lu0=-8.5946913e-011 pu0=1.9138983e-017             lvsat=0.0022891141               pvsat=-9.3503764e-011 lpclm=-5.4593543e-008            ppclm=4.8619973e-015             lbigc=1.6049542e-010 pbigc=-2.4200256e-017            lbigsd=3.4356646e-011             pbigsd=-3.363821e-018 lute=-2.0511044e-008            pute=6.2096135e-015             lat=-0.0004895385 pat=-4.009667e-011             leta0=0                          peta0=0 letab=1.5113261e-009             petab=-7.3052912e-017 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.005                      lvoff_mcl=-4.9e-16                   wvoff_mcl=-5.4e-15 pvoff_mcl=-1.7e-22                   ua1_ff=8.13992e-11                lua1_ff=-4.06996e-18 wua1_ff=-9.27951e-18               pua1_ff=4.63975e-25 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.27 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.63653423 lvth0=-3.7275135e-009            wvth0=-1.573974e-008             pvth0=1.0070452e-015 k2=-0.029418682               lk2=-1.8403028e-009            wk2=-4.0250586e-009 pk2=2.672288e-016              cit=0.013524026                voff=-0.28422312 lvoff=2.0294023e-009             wvoff=1.3667925e-008             pvoff=-6.1489202e-016 eta0=-0.0058600823              weta0=8.2004938e-010             etab=0.004640535 wetab=-4.338331e-009             u0=0.043520745                wu0=-3.9080176e-009 ua=-1.3105625e-009            lua=8.3395119e-018             wua=-1.5307126e-016 pua=9.8239197e-024             ub=2.0449829e-018             lub=-4.0469109e-026 wub=4.905298e-026              pub=-6.3036872e-033            uc=-4.0604315e-010 luc=1.4355491e-017             wuc=4.4164593e-017             puc=-2.2257096e-024 vsat=175912.45                  wvsat=-0.009925768               a0=7.2863172 la0=-6.9264539e-007            wa0=2.4188177e-008             pa0=-1.1091552e-014 ags=2.8518519                  lags=0                          wags=-9.7111111e-008 pags=0                          keta=-0.98566258                lketa=3.5986833e-008 wketa=1.6125887e-007             pketa=-8.2571656e-015            pclm=1.8722222 wpclm=-1.1653333e-007            pdiblc2=0.0023518519               wpdiblc2=-9.7111111e-011 aigbacc=0.0092259358               laigbacc=-6.6901608e-011            waigbacc=-1.4863324e-010 paigbacc=8.1843604e-018             aigc=0.012913586                laigc=-1.0263129e-010 waigc=-3.5021898e-010            paigc=8.9059417e-018             bigc=0.0049679019 wbigc=-4.4498918e-010            aigsd=0.0094759977               laigsd=2.4664631e-012 waigsd=-1.7630675e-011            paigsd=6.7307223e-019             bigsd=0.0014631276 wbigsd=-1.6797201e-010            tvoff=0.00290237                 ltvoff=-3.34051e-011 wtvoff=-2.26569e-010              ptvoff=1.09074e-017               kt1=-0.0092306724 lkt1=6.7030437e-010             wkt1=-2.0961188e-008            pkt1=8.8799067e-016 kt2=-0.052842145               lkt2=3.197668e-010              wkt2=2.8881417e-010 pkt2=8.2203484e-017             ute=-0.11399177                wute=-1.5483827e-007 ua1=-8.8435283e-010            lua1=-7.3253823e-017            wua1=3.7010183e-016 pua1=-1.3516628e-023            ub1=2.6419542e-018             lub1=2.2349326e-026 wub1=-7.7873056e-025            pub1=3.3192406e-032             uc1=1.0243489e-009 luc1=-2.2995221e-017            wuc1=-1.1728244e-016            puc1=4.6987885e-024 at=31453.743                  wat=0.006969402                lcit=-3.9981243e-010 wcit=-1.4724979e-009            pcit=6.6341564e-017             lu0=-1.1274873e-009 pu0=1.9776068e-016             lvsat=-0.0022672122              pvsat=5.574472e-010 lpclm=-6.9851852e-008            ppclm=7.9631111e-015             lbigc=-1.2620078e-010 pbigc=1.3079548e-017             lbigsd=-3.4887119e-011            pbigsd=7.4410849e-018 lute=-2.8050412e-008            pute=7.7419136e-015             lat=-0.00036311311 pat=-2.6886381e-010            leta0=2.2355967e-009             peta0=-1.7695802e-016 letab=-1.018386e-009             petab=2.0560311e-016 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' voff_mcl=0.00500001                 lvoff_mcl=-3.3e-16                   wvoff_mcl=-6e-16 pvoff_mcl=5.3e-22                    ua1_fs=-9.11108e-11               lua1_fs=4.55556e-18 wua1_fs=-2e-24                     pua1_fs=1.2e-31 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_hvt_mac.28 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.43024324 lvth0=4.7304176e-009             wvth0=1.7960492e-008             pvth0=-3.7466427e-016 k2=-0.078888313               lk2=1.8795207e-010             wk2=2.3068781e-009 pk2=7.6193963e-018             cit=-0.010099746               voff=-0.12398488 lvoff=-4.5403655e-009            wvoff=-1.4324375e-008            pvoff=5.3279227e-016 eta0=0.051958848                weta0=-8.3299753e-009            etab=-0.054931274 wetab=3.0561779e-009             u0=0.0019693044               wu0=3.3891853e-009 ua=-3.3576688e-009            lua=9.2270872e-017             wua=2.8264633e-016 pua=-8.0405015e-024            ub=3.268969e-018              lub=-9.0652537e-026 wub=-3.144045e-025             pub=8.5980694e-033             uc=5.2644634e-011 luc=-4.4507083e-018            wuc=-2.2613695e-017            puc=5.1220016e-025 vsat=-14093.306                 wvsat=0.013287685                a0=-9.4488382 la0=-6.5040213e-009            wa0=3.2149216e-008             pa0=-1.1417955e-014 ags=2.8518519                  lags=0                          wags=-9.7111111e-008 pags=0                          keta=0.48867677                 lketa=-2.446108e-008 wketa=-9.5728117e-008            pketa=2.2793008e-015             pclm=0.0069303704 wpclm=2.379766e-007              pdiblc2=0.0023518519               wpdiblc2=-9.7111111e-011 aigbacc=0.0062552799               laigbacc=5.4895281e-011             waigbacc=2.8097704e-010 paigbacc=-9.4296611e-018            aigc=0.011722334                laigc=-5.3789943e-011 waigc=-1.3192443e-010            paigc=-4.413503e-020             bigc=0.0028327201 wbigc=-1.4814088e-010            aigsd=0.0088784002               laigsd=2.6967959e-011 waigsd=1.1597667e-010             paigsd=-4.8048288e-018            bigsd=-0.00013552428 wbigsd=1.857455e-010              tvoff=0.0020242                  ltvoff=2.5997e-012 wtvoff=1.70605e-010               ptvoff=-5.37669e-018              kt1=-0.090859772 lkt1=4.0170975e-009             wkt1=1.4227033e-008             pkt1=-5.5472641e-016 kt2=-0.097284611               lkt2=2.1419079e-009             wkt2=5.443567e-009 pkt2=-1.2914138e-016            ute=0.12695473                 wute=-5.3950617e-010 ua1=1.7687119e-009             lua1=-1.8202948e-016            wua1=-2.4301262e-016 pua1=1.1621065e-023             ub1=-6.8686122e-019            lub1=1.5883076e-025 wub1=2.821993e-025              pub1=-1.0305718e-032            uc1=5.6769591e-010 luc1=-4.2724497e-018            wuc1=4.6506133e-017             puc1=-2.0165429e-024 at=35316.932                  wat=-0.004674257               lcit=5.6876226e-010 wcit=1.4228634e-009             pcit=-5.236825e-017             lu0=5.7612181e-010 pu0=-1.0142464e-016            lvsat=0.0055230237               pvsat=-3.9430438e-010 lpclm=6.6251141e-009             ppclm=-6.5717963e-015            lbigc=-3.8658326e-011 pbigc=9.0876794e-019             lbigsd=3.0657607e-011             pbigsd=-7.061333e-018 lute=-3.7929218e-008            pute=1.4156642e-015             lat=-0.00052150385 pat=2.0852621e-010             leta0=-1.3497942e-010            peta0=1.9819299e-016 letab=1.4240581e-009             petab=-9.7571758e-017 jtsswgs='7.6e-006*(1+0.645*iboffn_flag_hvt)'                               jtsswgd='7.6e-006*(1+0.645*iboffn_flag_hvt)' vth0_mc=0.0302881                  lvth0_mc=-1.24181e-09               wvth0_mc=-3.45284e-09 pvth0_mc=1.41566e-16                voff_ff=-0.0121152                 voff_mcl=0.0175103 voff_mc=0.0302881                  lvoff_ff=4.96724e-10                lvoff_mcl=-5.12921e-10 lvoff_mc=-1.24181e-09               wvoff_ff=1.38114e-09                wvoff_mcl=-3.45284e-09 wvoff_mc=-3.45284e-09               pvoff_ff=-5.66266e-17               pvoff_mcl=1.41566e-16 pvoff_mc=1.41566e-16                u0_mc=-0.00658436                wu0_mc=3.45282e-10 ua_ff=-1.21152e-10               lua_ff=4.96724e-18                wua_ff=1.38114e-17 pua_ff=-5.66266e-25               vsat_ff=1251.03                    vsat_fs=-6057.61 vsat_mc=50567.9                    wvsat_ff=-0.000345284               wvsat_fs=0.000690568 wvsat_mc=-0.00414341                ua1_fs=9.11108e-11                lua1_fs=-2.91555e-18 wua1_fs=2e-24                      pua1_fs=3.2e-31                    lu0_mc=2.69959e-10 pu0_mc=-1.41566e-17               lvsat_ff=-5.12922e-05               lvsat_fs=0.000248362 lvsat_mc=-0.00207328                pvsat_ff=1.41566e-11                pvsat_fs=-2.83133e-11 pvsat_mc=1.6988e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model pch_hvt_mac.global pmos ( modelid=4                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_hvt'             permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=2.18e-009                  toxm=2.18e-009                  dtox=4.69e-010 epsrox=3.9                        wint=0                          lint=0 ll=0                          wl=0                          lln=1 wln=1                          lw=0                          ww=0 lwn=1                          wwn=1                          lwl=0 wwl=0                          llc=0                          wlc=0 lwc=0                          wwc=0                          lwlc=0 wwlc=0                          xl=-3e-009                    xw=6e-009 dlc=5.66905e-009               dwc=0                          xpart=1 toxref=3e-009                     dlcig=2.5e-009                   k1=0.46526 k3=-2.835                     k3b=1.5                        w0=0 dvt0=4                          dvt1=1.85                       dvt2=0.03 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.4492                    voffl=0 dvtp0=6.2688e-007                dvtp1=0.015                      lpe0=0 lpeb=-8.909e-009                xj=8.5e-008                   ngate=1.1e+020 ndep=6e+017                     nsd=1e+020                     phin=0.1615 cdsc=0                          cdscb=0                          cdscd=0 nfactor=1                          ud=0                          lud=0 wud=0                          pud=0                          a1=0 a2=1                          b0=0                          b1=0 dwg=0                          dwb=0                          pdiblc1=0 pdiblcb=0                          drout=0.56                       pvag=0.03 delta=0.018814                   pscbe1=9.264e+008                 pscbe2=1e-020 fprout=200                        pdits=0                          pditsd=0 pditsl=0                          rsh=16.7                       rdsw=160 rsw=100                        rdw=100                        prwg=0 prwb=0                          wr=1                          alpha0=4.4e-006 alpha1=2                          beta0=19.2                       agidl=3.5e-010 bgidl=1.38e+009                  cgidl=0.2                        egidl=0.001 bigbacc=0.006                      cigbacc=0.245                      nigbacc=10 bigbinv=0.00149                    cigbinv=0.006                      eigbinv=1.1 nigbinv=2.1927                     cigc=0.15259                    cigsd=0.0011 nigc=2.291                      poxedge=1                          pigcd=3.15 ntox=1                          xrcrg1=12                         xrcrg2=1 vfbsdoff=0.01                       lvfbsdoff=0                          wvfbsdoff=0 pvfbsdoff=0                          cgso=4.92779e-011               cgdo=4.92779e-011 cgbo=0                          cgdl=4.63343e-011               cgsl=4.63343e-011 clc=0                          cle=0.6                        cf='9e-11+0.92e-10*ccoflag_hvt' ckappas=0.6                        ckappad=0.6                        acde=0.4 moin=8.731                      noff=2.3488                     voffcv=-0.084 tvfbsdoff=0.114                      ltvfbsdoff=0                          wtvfbsdoff=0 ptvfbsdoff=0                          kt1l=0                          prt=0 fnoimod=1                          tnoimod=0                          em=2e+007 ef=1.18                       noia=0                          noib=0 noic=0                          lintnoi=-2.17e-008                 jss=8.95e-07 jsd=8.95e-07                   jsws=2.11e-13                   jswd=2.11e-13 jswgs=2.11e-13                   jswgd=2.11e-13                   njs=1.02 njd=1.02                       ijthsfwd=0.01                       ijthdfwd=0.01 ijthsrev=0.01                       ijthdrev=0.01                       bvs=7.000000e+00 bvd=7.000000e+00               xjbvs=1                          xjbvd=1 njtsswg=10                         xtsswgs=0.13                       xtsswgd=0.13 tnjtsswg=1                          vtsswgs=0.77008                    vtsswgd=0.77008 pbs=0.938                      pbd=0.938                      cjs=0.001739 cjd=0.001739                   mjs=0.518                      mjd=0.518 pbsws=0.777                      pbswd=0.777                      cjsws=1.242e-010 cjswd=1.242e-010                 mjsws=0.253                      mjswd=0.253 pbswgs=0.907                      pbswgd=0.907                      cjswgs=3e-010 cjswgd=3e-010                     mjswgs=0.6                        mjswgd=0.6 tpb=0.00096                    tcj=0.00069                    tpbsw=0.00061 tcjsw=0.00021                    tpbswg=0.00062                    tcjswg=0.00075 xtis=3                          xtid=3                          dmcg=3.75e-008 dmci=3.75e-008                  dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=-5.10e-009 rshg=14.4                       gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          lnfactor=0 pnfactor=0                          wnfactor=0                          k2we=0 ku0we=-0.0004                    kvth0we=-0.0004346                 lk2we=0e-11 lku0we=-1e-11                     lkvth0we=1e-011                     pk2we=0e-18 pku0we=2e-18                      pkvth0we=-1.063e-019                scref=1e-6 web=2251.7                     wec=-7896.1                    wk2we=0e-11 wku0we=-1e-010                    wkvth0we=-7e-012                    wpemod=1 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.2                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.6 bidirectionflag='bidirectionflag_mos_hvt' iboffn_flag='iboffn_flag_hvt' iboffp_flag='iboffp_flag_hvt' sigma_factor='sigma_factor_hvt' ccoflag='ccoflag_hvt' rcoflag='rcoflag_hvt' rgflag='rgflag_hvt' mismatchflag='mismatchflag_mos_hvt' globalflag='globalflag_mos_hvt' totalflag='totalflag_mos_hvt' designflag='designflag_mos_hvt' global_factor='global_factor_hvt' local_factor='local_factor_hvt' sigma_factor_flicker='sigma_factor_flicker_hvt' noiseflag='noiseflagp_hvt' noiseflag_mc='noiseflagp_hvt_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w31='2.3875*0.35355' w32='0.70711*0.35355' w33='0.54772*0.31715' w34='0.54772*0.2225' w35='0.54772*-0.17742' w36='0.54772*-0.6346' w37='0.54772*0.40656' w38='0.54772*0.020451' w39='0' w40='0' tox_c='toxp_hvt'                 ntox_c='ntoxp_hvt'                dxl_c='dxlp_hvt' dxw_c='dxwp_hvt'                 cj_c='cjp_hvt'                  cjsw_c='cjswp_hvt' cjswg_c='cjswgp_hvt'               cgo_c='cgop_hvt'                 cgl_c='cglp_hvt' ddlc_c='ddlcp_hvt'                dvth_c='dvthp_hvt'                dlvth_c='dlvthp_hvt' dwvth_c='dwvthp_hvt'               dpvth_c='dpvthp_hvt'               dk2_c='dk2p_hvt' dlk2_c='dlk2p_hvt'                dwk2_c='dwk2p_hvt'                dpk2_c='dpk2p_hvt' deta0_c='deta0p_hvt'               dleta0_c='dleta0p_hvt'              dweta0_c='dweta0p_hvt' dpeta0_c='dpeta0p_hvt'              dvoff_c='dvoffp_hvt'               dlvoff_c='dlvoffp_hvt' dwvoff_c='dwvoffp_hvt'              dpvoff_c='dpvoffp_hvt'              dcit_c='dcitp_hvt' dlcit_c='dlcitp_hvt'               dwcit_c='dwcitp_hvt'               dpcit_c='dpcitp_hvt' dnfactor_c='dnfactorp_hvt'            dlnfactor_c='dlnfactorp_hvt'           dwnfactor_c='dwnfactorp_hvt' dpnfactor_c='dpnfactorp_hvt'           du0_c='du0p_hvt'                 dlu0_c='dlu0p_hvt' dwu0_c='dwu0p_hvt'                dpu0_c='dpu0p_hvt'                dub_c='dubp_hvt' dlub_c='dlubp_hvt'                dwub_c='dwubp_hvt'                dpub_c='dpubp_hvt' dpclm_c='dpclmp_hvt'               dlpclm_c='dlpclmp_hvt'              dwpclm_c='dwpclmp_hvt' dppclm_c='dppclmp_hvt'              dvsat_c='dvsatp_hvt'               dlvsat_c='dlvsatp_hvt' dwvsat_c='dwvsatp_hvt'              dpvsat_c='dpvsatp_hvt'              da0_c='da0p_hvt' dla0_c='dla0p_hvt'                dwa0_c='dwa0p_hvt'                dpa0_c='dpa0p_hvt' dags_c='dagsp_hvt'                dlags_c='dlagsp_hvt'               dwags_c='dwagsp_hvt' dpags_c='dpagsp_hvt'               dpkt1_c='dpkt1p_hvt'               dat_c='datp_hvt' dlat_c='dlatp_hvt'                dwat_c='dwatp_hvt'                dpat_c='dpatp_hvt' dua1_c='dua1p_hvt'                dlua1_c='dlua1p_hvt'               dwua1_c='dwua1p_hvt' dpua1_c='dpua1p_hvt'               cf_c='cfp_hvt'                  jtsswg_c='jtsswgp_hvt' dpdiblc2_c='dpdiblc2p_hvt'            dminv_c='dminvp_hvt'               dketa_c='dketap_hvt' dlketa_c='dlketap_hvt'              dwketa_c='dwketap_hvt'              dpketa_c='dpketap_hvt' ss_flag_c='ss_flagp_hvt'             ff_flag_c='ff_flagp_hvt'             sf_flag_c='sf_flagp_hvt' fs_flag_c='fs_flagp_hvt'             monte_flag_c='monte_flagp_hvt'         c1f_c='c1fp_hvt' c2f_c='c2fp_hvt'                 c3f_c='c3fp_hvt' global_mc='global_mc_flag_hvt' tox_g='toxp_hvt_ms_global'       ntox_g='ntoxp_hvt_ms_global'      dxl_g='dxlp_hvt_ms_global' dxw_g='dxwp_hvt_ms_global'       cj_g='cjp_hvt_ms_global'        cjsw_g='cjswp_hvt_ms_global' cjswg_g='cjswgp_hvt_ms_global'     cgo_g='cgop_hvt_ms_global'       cgl_g='cglp_hvt_ms_global' dvth_g='dvthp_hvt_ms_global'      dlvth_g='dlvthp_hvt_ms_global' dwvth_g='dwvthp_hvt_ms_global'     dpvth_g='dpvthp_hvt_ms_global'     dk2_g='dk2p_hvt_ms_global' dleta0_g='dleta0p_hvt_ms_global'    du0_g='du0p_hvt_ms_global'       dlu0_g='dlu0p_hvt_ms_global' dwu0_g='dwu0p_hvt_ms_global'      dpu0_g='dpu0p_hvt_ms_global' dpclm_g='dpclmp_hvt_ms_global'     dvsat_g='dvsatp_hvt_ms_global' dlvsat_g='dlvsatp_hvt_ms_global'    dwvsat_g='dwvsatp_hvt_ms_global' dpvsat_g='dpvsatp_hvt_ms_global'    dags_g='dagsp_hvt_ms_global' dwags_g='dwagsp_hvt_ms_global'     dpkt1_g='dpkt1p_hvt_ms_global'     dat_g='datp_hvt_ms_global' dua1_g='dua1p_hvt_ms_global'      dlua1_g='dlua1p_hvt_ms_global' dpua1_g='dpua1p_hvt_ms_global'     cf_g='cfp_hvt_ms_global' dpdiblc2_g='dpdiblc2p_hvt_ms_global'  dminv_g='dminvp_hvt_ms_global' dlketa_g='dlketap_hvt_ms_global'    ss_flag_g='ss_flagp_hvt_ms_global' ff_flag_g='ff_flagp_hvt_ms_global'   monte_flag_g='monte_flagp_hvt_ms_global' sf_flag_g='sf_flagp_hvt_ms_global'   fs_flag_g='fs_flagp_hvt_ms_global' weight1=-3.2636667 weight2=2.053 weight3=1.1308667 weight4=0.66666667 weight5=-0.46406 tox_1=4.3294216e-012 tox_2=-1.000905e-011 tox_3=-8.7172436e-013 tox_4=-3.7477187e-011 tox_5=7.390037e-013 ntox_1=0.020071 ntox_2=-0.0059138 ntox_3=-0.0019932 ntox_4=9.2745e-018 ntox_5=-0.0017413 dxl_1=9.802549e-011 dxl_2=-2.2662113e-010 dxl_3=-1.9737099e-011 dxl_4=8.4853424e-010 dxl_5=1.6732084e-011 dxw_1=-7.2934365e-010 dxw_2=-8.2157411e-010 dxw_3=2.5306127e-011 dxw_4=-1.2950065e-024 dxw_5=-5.8959295e-009 dxw_max=-3.5e-008 cj_1=1.2216e-005 cj_2=-3.5994e-006 cj_3=-1.2132e-006 cj_4=-1.0385e-020 cj_5=-1.0598e-006 cjsw_1=8.7248e-013 cjsw_2=-2.5707e-013 cjsw_3=-8.6646e-014 cjsw_4=2.127e-029 cjsw_5=-7.5693e-014 cjswg_1=2.1074e-012 cjswg_2=-6.2095e-013 cjswg_3=-2.0929e-013 cjswg_4=-1.4206e-028 cjswg_5=-1.8283e-013 cgo_1=-3.4617e-013 cgo_2=1.02e-013 cgo_3=3.4378e-014 cgo_4=-3.9359e-028 cgo_5=3.0032e-014 cgl_1=-3.2549e-013 cgl_2=9.5904e-014 cgl_3=3.2324e-014 cgl_4=2.6329e-028 cgl_5=2.8238e-014 dvth_1=-0.0027678 dvth_2=-0.0041278 dvth_3=2.4813e-005 dvth_4=-1.8436e-018 dvth_5=0.00087104 dlvth_1=-1.4397e-010 dlvth_2=1.3294e-012 dlvth_3=3.1814e-011 dlvth_4=1.6837e-025 dlvth_5=1.6412e-011 dwvth_1=-1.4617e-010 dwvth_2=4.391e-011 dwvth_3=-5.0467e-011 dwvth_4=-2.0436e-026 dwvth_5=1.2117e-011 dpvth_1=-2.657e-017 dpvth_2=-2.472055e-017 dpvth_3=1.9859e-018 dpvth_4=-2.7938e-032 dpvth_5=6.2946e-018 dk2_1=0.00063244 dk2_2=0.0009671 dk2_3=-4.4609e-006 dk2_4=-9.2167e-020 dk2_5=-0.00020208 dleta0_1=-4.0142e-011 dleta0_2=1.1828e-011 dleta0_3=3.9865e-012 dleta0_4=8.3187e-027 dleta0_5=3.4826e-012 du0_1=5.7263e-005 du0_2=0.00014796 du0_3=-1.2506e-006 du0_4=-1.726e-020 du0_5=-2.6032e-005 dlu0_1=3.2677e-013 dlu0_2=1.5584e-012 dlu0_3=-4.8196e-013 dlu0_4=6.689e-028 dlu0_5=-2.4328e-013 dwu0_1=8.6648e-012 dwu0_2=6.5303e-012 dwu0_3=7.7821e-013 dwu0_4=-1.1874e-026 dwu0_5=-2.0487e-012 dpu0_1=-8.3423e-020 dpu0_2=2.3714e-018 dpu0_3=3.5862e-019 dpu0_4=-1.0585e-033 dpu0_5=-4.6587e-019 dpclm_1=-0.0050177 dpclm_2=0.0014784 dpclm_3=0.00049831 dpclm_4=-4.6809e-018 dpclm_5=0.00043532 dvsat_1=167.34 dvsat_2=1427.6 dvsat_3=-21.698 dvsat_4=6.7386e-013 dvsat_5=-174.37 dlvsat_1=3.0267e-005 dlvsat_2=-8.8088e-006 dlvsat_3=-1.1441e-005 dlvsat_4=-2.9206e-020 dlvsat_5=-2.6991e-006 dwvsat_1=3.0264e-005 dwvsat_2=0.0002584 dwvsat_3=5.8389e-005 dwvsat_4=-1.7542e-019 dwvsat_5=-5.3928e-005 dpvsat_1=3.6001e-012 dpvsat_2=-1.0318e-012 dpvsat_3=-2.5929e-012 dpvsat_4=2.1248e-027 dpvsat_5=-3.3175e-013 dags_1=0.052626 dags_2=0.050405 dags_3=-0.0018922 dags_4=2.5496e-017 dags_5=-0.012978 dwags_1=2.4267e-010 dwags_2=2.0706e-009 dwags_3=8.4258e-011 dwags_4=1.2201e-025 dwags_5=-2.9445e-010 dpkt1_1=2.5748e-018 dpkt1_2=-8.4275e-019 dpkt1_3=6.2426e-018 dpkt1_4=-2.7551e-033 dpkt1_5=-1.6694e-019 dat_1=1089.8 dat_2=-309.49 dat_3=-1005 dat_4=-1.0994e-012 dat_5=-102.33 dua1_1=1.0035e-011 dua1_2=-2.9569e-012 dua1_3=-9.9661e-013 dua1_4=5.6481e-027 dua1_5=-8.7064e-013 dlua1_1=-7.8954e-020 dlua1_2=3.4364e-020 dlua1_3=-8.4994e-019 dlua1_4=8.2293e-035 dlua1_5=-6.0046e-022 dpua1_1=-8.0283e-026 dpua1_2=2.3655e-026 dpua1_3=7.9729e-027 dpua1_4=-1.0198e-041 dpua1_5=6.9651e-027 cf_1=-6.3223e-013 cf_2=1.8628e-013 cf_3=6.2787e-014 cf_4=-7.0189e-029 cf_5=5.485e-014 dpdiblc2_1=-2.0071e-005 dpdiblc2_2=5.9138e-006 dpdiblc2_3=1.9932e-006 dpdiblc2_4=5.2331e-021 dpdiblc2_5=1.7413e-006 dminv_1=-0.011501 dminv_2=0.0033383 dminv_3=0.0050412 dminv_4=-4.0506e-018 dminv_5=0.0010317 dlketa_1=-5.1496e-010 dlketa_2=1.6855e-010 dlketa_3=-1.2485e-009 dlketa_4=-2.6853e-025 dlketa_5=3.3388e-011 ss_flag_1=0.048858 ss_flag_2=-0.012714 ss_flag_3=-0.13482 ss_flag_4=6.157e-017 ss_flag_5=-0.0053676 ff_flag_1=-0.051496 ff_flag_2=0.016855 ff_flag_3=-0.12485 ff_flag_4=1.8969e-017 ff_flag_5=0.0033388 monte_flag_1=0.0816875 monte_flag_2=-0.18885 monte_flag_3=-0.0164475 monte_flag_4=0.707108 monte_flag_5=0.0139433 sigma_local=1                          a_1=0.918491 b_1=-7.32652e-005              c_1=0.00235899                 d_1=0.000085966 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1.0575                     b_2=-0.00482861                c_2=-0.00257128 d_2=-0.000454853               a_3=0.976279                   b_3=-0.00672237 c_3=-0.00200969                d_3=-0.000232988               e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.85 b_4=-0.001                     c_4=-0.01                      d_4=-0.0003 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=0.84                       b_5=-0.004                     c_5=-0.01 d_5=-0.0003                    e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=-0.0016                    mis_a_2=-0.071                     mis_a_3=0.039 mis_b_1=0.002                      mis_b_2=-0.2                       mis_b_3=0.0212 mis_c_1=0.1                        mis_c_2=0                          mis_c_3=0 mis_d_1=0.00076                    mis_d_2=0                          mis_d_3=0 mis_e_1=0.0018                     mis_e_2=0.287                      mis_e_3=-0.131 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-3e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=60                         co_rsd=16.7 cf0=9e-11                      cco=0.92e-10 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.5                        l_rjtsswg=0.005                      ll_rjtsswg=1 w_rjtsswg=0.5                        ww_rjtsswg=1.0                        p_rjtsswg=0.0 noimod=1                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6               sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=1                   lreflod=0.9e-6              llodref=2 lod_clamp=-1e90 wlod0=0 ku00=-0e-9       lku00=0e-7        wku00=0e-8         pku00=0e-14 tku00=0           llodku00=1           wlodku00=1            kvsat0=0.5 kvth00=-3.8e-9     lkvth00=1.75e-8     wkvth00=3e-8         pkvth00=0e-15 llodvth0=1           wlodvth0=1 stk20=0           lodk20=1           steta00=5e-11        lodeta00=1 wlod00=0 ku000=0           lku000=-13e-32     wku000=0            pku000=0 llodku000=3           wlodku000=1 kvth000=0           lkvth000=3e-17       wkvth000=0            pkvth000=0e-14 llodvth00=1           wlodvth00=1 steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0           llod1=0.00e-6 ku01=2e-8        lku01=-3e-2       wku01=-5e-15     pku01=0 llodku01=-1          wlodku01=1           kvsat1=-0 kvth01=11e-9     lkvth01=-3e-24      wkvth01='1.5e-19'     pkvth01=0e-24 llodvth1=2           wlodvth1=1.5 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.1        lku02=0.4e-7      wku02=0            pku02=0 tku02=0           llodku02=1           wlodku02=1            kvsat2='0.4*0+0.5' kvth02=-0e-3       lkvth02=0e-8        wkvth02=0e-8         pkvth02=0 llodvth2=1           wlodvth2=1 stk22=0           lodk22=1           steta02=-1e-4        lodeta02=1 wlod02=0 ku002=0           lku002='-1.2e11*2'     wku002=3.5e-9       pku002=0 llodku002=-2          wlodku002=1 kvth002=0           lkvth002=-0e-11      wkvth002=0            pkvth002=0 llodvth02=1           wlodvth02=1 steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0.085        lku03=-0.05e-7        wku03=0e-7         pku03=0 tku03=0           llodku03=1           wlodku03=1            kvsat3=0.4 kvth03=0.1e-3      lkvth03=0e-20       wkvth03=0e-8         pkvth03=0e-20 llodvth3=3           wlodvth3=1 stk23=0           lodk23=1           steta03=0e-3         lodeta03=1 wlod03=0 ku003=0           lku003='-1.25e5*8e-1'     wku003=1.5e-9            pku003=0 llodku003=-1          wlodku003=1 kvth003=0e-3        lkvth003=-5e-26      wkvth003=-2e-10       pkvth003=0e-32 llodvth03=3           wlodvth03=1 steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.7                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=-1.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=-0.000              wkvth0dpl=0                   wdplkvth0=1 lkvth0dpl=0.0e-9              ldplkvth0=1.0                 pkvth0dpl=0 ku0dpl=1               wku0dpl=0                   wdplku0=1 lku0dpl=-4e-8              ldplku0=1                 pku0dpl=0 keta0dpl=0.00                wketa0dpl=0                   wdplketa0=1 kvsatdpl=0                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=1 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=1.0e-6              wkvth0dpx=0                   wdpxkvth0=1 lkvth0dpx=0                   ldpxkvth0=1                   pkvth0dpx=0 ku0dpx=0                   wku0dpx=0                   wdpxku0=1 lku0dpx=0                   ldpxku0=1                   pku0dpx=0 keta0dpx=0                   wketa0dpx=0                   wdpxketa0=1 kvsatdpx=0                   wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0.02               wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-2             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='0.5'               wku0dps=0                   wdpsku0=1 lku0dps='2e-8+0e-8'        ldpsku0=1.0                 pku0dps=0 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0.7                 wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=1 ku0dps_b1=0                 ku0dps_b2=0.11 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=0.002               wkvth0dpa=-2.0e-9            wdpakvth0=1 lkvth0dpa=0.015e-7            ldpakvth0=1.0                pkvth0dpa=-3.0e-17 ku0dpa=-0.1               wku0dpa=2e-9               wdpaku0=1 lku0dpa=-7e-9               ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=1 ku0dpa_b1=-0.1             ku0dpa_b2=0.00 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2=-0.01               wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0.5e-9              ldp2kvth0=1                   pkvth0dp2=0 ku0dp2=0.1                wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=-0.0e-8              ldp2ku0=1.0                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0.00                wdp2=0 kvth0dp2l=-0.018              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.6               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0e-8               ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0.2                wdp2l=0 kvth0dp2l_b1=0.00            kvth0dp2l_b2=-0.016           dp2lbinflg=1 ku0dp2l_b1=-0.00            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=-0.007              wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=-0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.2              wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=-25.0e-5            ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=0.017           kvth0dp2a_b2=-0.02           dp2abinflg=1 ku0dp2a_b1=-0.12                ku0dp2a_b2=0.08 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx=-0.023              wkvth0enx=-0.0e-9             wenxkvth0=1.0 lkvth0enx=-11.0e-9              lenxkvth0=1.0                 pkvth0enx=-0.85e-16 ku0enx=-2.0                wku0enx=-1.0e-8             wenxku0=1.0 lku0enx=0.4e-7              lenxku0=1.0                 pku0enx=-7.0e-16 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=1.0                 wka0enx=0                   wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx=0.5                 wenx=0                   ku0enx0=-0.20 eny0=0.08e-6 enyref=0.08e-6             enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0.010               wkvth0eny=5.0e-10             wenykvth0=1 lkvth0eny=1.0e-8              lenykvth0=1.0                 pkvth0eny=0 ku0eny=14.0                wku0eny=1.0e-8              wenyku0=1 ku0eny0=0.04                wku0eny0=-1.0e-7             weny0ku0=1 lku0eny=8.0e-6              lenyku0=1.0                 pku0eny=2.0e-16 keta0eny=0e-4                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny=0.8                 weny=0 kvth0eny1=-6e-4              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=3.0e-18 ku0eny1=-1.5e-3            wku0eny1=-1.0e-10           weny1ku0=1 lku0eny1=-0.6e-8            leny1ku0=1.0                pku0eny1=-5.5e-17 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1=1.0e-8             weny1ka0=1 lka0eny1=4.0e-9             leny1ka0=1.0                pka0eny1=1.5e-15 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=0.045               wkvth0rx=0.0e-6              wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0e-15 ku0rx=0.05                wku0rx=0.0e-4              wrxku0=1.0 lku0rx=0.0e-7              lrxku0=1.0                 pku0rx=0.0e-14 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.4                 wrx=0                   ku0rx0=0.35 ry_mode=0 ryref=1.8027e-5           ringymax=1.8047e-5           ringymin=0.117e-6 kvth0ry=-0.0025             wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry='1.0e-8*0'           lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry=-0.8                 wku0ry=-0.5e-8             wryku0=1.0 lku0ry=4.0e-7               lryku0=1.0                 pku0ry=-2.0e-16 keta0ry=0.00                 wketa0ry=0                   wryketa0=1 kvsatry=0.7                 wry=0 kvth0ry0='-0.01*0'            ku0ry0='-0.14*0' sfxref=9.0e-8            sfxmax=1.53e-6          minwodx=0 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=0.0 kvth0odx1a=-0.009            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.1               lku0odx1a=1.6e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.6 kvth0odx1b=0.0000            lkvth0odx1b=2.7e-11           lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.0004           lku0odx1b=1.25e-6           lodx1bku0=0.5 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6 sfymax=1.53e-6           minwody=0.0e-6            wody=5e-7 kvth0odya=50                lkvth0odya=1.0e-4            lodyakvth0=1.0 wkvth0odya=1.8e-7            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=1.5                 lku0odya=1.0e-6            lodyaku0=1.0 wku0odya=-0.0e-8           wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=-11e-2           wketa0ody=0                 wodyketa0=1 kvsatody=0 lrefody=1.0e-7            lodyref=1 kvth0odyb=-0.00             lkvth0odyb=7.0e-17           lodybkvth0=2.0 wkvth0odyb=9.0e-9            wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.55             lku0odyb=4.5e-10           lodybku0=1.1 wku0odyb=-0.9e-7           wodybku0=1.0               pku0odyb=-1.8e-16 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model pch_hvt_mac.1 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.46206573 lvth0=1.286056e-008              wvth0=-2.9750667e-008            pvth0=1.1502568e-014 k2=0.027255346                lk2=2.7235547e-009             wk2=-2.2032688e-008 pk2=2.9114425e-015             cit=0.0022371275               lcit=7.6825057e-014 wcit=-7.8135562e-010            pcit=-1.0256934e-019            voff=-0.13182743 lvoff=1.019023e-011              wvoff=-1.334748e-008             pvoff=-1.1265181e-017 eta0=0.12                       etab=-0.05469247                wetab=-6.8228622e-008 u0=0.0097467                  wu0=2.956278e-010              ua=3.600425e-010 lua=-3.7649312e-016            wua=-4.1622152e-016            pua=1.669774e-022 ub=8.5908199e-019             lub=4.8540667e-026             wub=3.8084506e-025 pub=-2.5166465e-032            uc=-5.4810135e-010            luc=4.3276783e-016 wuc=9.0659192e-018             puc=-8.1566075e-023            vsat=87550 wvsat=-0.0113703                 a0=2.8253074                  la0=-7.2054907e-012 wa0=-1.0089103e-006            pa0=7.2503178e-018             ags=1.360535 lags=3.5427347e-007             wags=-4.5564578e-007            pags=1.443602e-013 keta=-0.47098473                lketa=3.1007921e-007             wketa=1.237914e-007 pketa=-4.9845935e-014            pclm=0.28109224                 lpclm=-4.0133298e-008 wpclm=-1.328667e-007             ppclm=3.6358674e-014             pdiblc2=0.0005 aigbacc=0.011409201                laigbacc=-4.1527772e-011            waigbacc=5.6397616e-010 paigbacc=-3.4177545e-017            aigbinv=0.00922051                 waigbinv=1.1347559e-009 aigc=0.0066563515               laigc=1.5641095e-011             waigc=-7.9211713e-010 paigc=9.4980069e-018             bigc=0.002173407                wbigc=-8.7710494e-010 aigsd=0.0047104825               laigsd=6.6792709e-012             waigsd=3.1061327e-010 paigsd=-6.0504355e-018            bigsd=4.095e-005                 wbigsd=2.387763e-010 tvoff=0.00290372                 ltvoff=-1.04137e-009              wtvoff=-2.34367e-011 ptvoff=-2.53575e-016              kt1=-0.33163924                lkt1=9.1846644e-008 wkt1=1.3607219e-007             pkt1=-1.2089827e-013            kt2=-0.06748513 wkt2=1.7653528e-008             ute=-1.6238665                 wute=6.0069295e-007 ua1=2.818326e-009              lua1=-1.112978e-015             wua1=-1.5966991e-016 pua1=1.0921538e-021             ub1=-3.2832044e-018            lub1=7.810465e-030 wub1=2.429843e-025              pub1=-8.8816393e-036            uc1=9.0707629e-012 luc1=5.6244059e-016             wuc1=1.5273389e-015             puc1=-2.1510375e-021 at=100000                     lu0=0                          pu0=0 lat=0                          wat=0                          pat=0 leta0=0                          weta0=0                          peta0=0 lvsat=0                          pvsat=0                          jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)' jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                ua1_ff=5.53018e-12 ua1_ss=-5.53018e-12               ua1_fs=-5.53018e-12               ua1_sf=5.53018e-12 lua1_ff=-4.98105e-17               lua1_ss=4.98105e-17                lua1_fs=4.98105e-17 lua1_sf=-4.98105e-17               wua1_ff=-3.2e-23                   wua1_ss=3.2e-23 wua1_fs=3.2e-23                    wua1_sf=-3.2e-23                   pua1_ff=7e-29 pua1_ss=-7e-29                     pua1_fs=-7e-29                     pua1_sf=7e-29 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.2 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.44123552 lvth0=-5.824148e-009             wvth0=-3.2834204e-008            pvth0=1.4268501e-014 k2=0.033954027                lk2=-3.2851623e-009            wk2=-1.6290663e-008 pk2=-2.2391542e-015            cit=0.00059415266              lcit=1.4738252e-009 wcit=3.939699e-010              pcit=-1.0543696e-015            voff=-0.12541642 lvoff=-5.7404888e-009            wvoff=-1.8245072e-008            pvoff=4.3818746e-015 eta0=0.12                       etab=-0.05469247                wetab=-6.8228622e-008 u0=0.0095162864               wu0=2.865922e-010              ua=3.8899765e-010 lua=-4.0246589e-016            wua=-3.5616918e-016            pua=1.1311046e-022 ub=6.4820483e-019             lub=2.3769748e-025             wub=6.2615898e-025 pub=-2.4521305e-031            uc=-1.2150507e-010            luc=5.0110965e-017 wuc=-2.765257e-017             puc=-4.8629591e-023            vsat=87550 wvsat=-0.0113703                 a0=3.9985914                  la0=-1.0524429e-006 wa0=-2.0766754e-006            pa0=9.5779261e-013             ags=1.9875329 lags=-2.0814363e-007            wags=-9.1985753e-007            pags=5.6075814e-013 keta=-0.1551                    lketa=2.67306e-008               wketa=6.82218e-008 pketa=9.9709614e-029             pclm=0.29507585                 lpclm=-5.2676594e-008 wpclm=-2.6060016e-007            ppclm=1.5093559e-013             pdiblc2=-0.0009146954 aigbacc=0.011305154                laigbacc=5.1802565e-011             waigbacc=1.0292132e-009 paigbacc=-4.5149515e-016            aigbinv=0.0091507791               waigbinv=9.2884414e-010 aigc=0.0079944166               laigc=-1.1846033e-009            waigc=-2.2871946e-009 paigc=1.3505825e-015             bigc=0.0037135842               wbigc=-2.6196201e-009 aigsd=0.0042466251               laigsd=4.2275937e-010             waigsd=7.9122897e-010 paigsd=-4.3716271e-016            bigsd=-0.00044453173             wbigsd=7.4476981e-010 tvoff=0.00201573                 ltvoff=-2.44844e-010              wtvoff=-7.72557e-010 ptvoff=4.18386e-016               kt1=-0.20551991                lkt1=-2.1282396e-008 wkt1=-2.6329839e-008            pkt1=2.4776347e-014             kt2=-0.07284099 wkt2=2.2375585e-008             ute=-2.351142                  wute=1.4887793e-006 ua1=9.5529866e-010             lua1=5.5815759e-016             wua1=3.7040096e-015 pua1=-2.3735667e-021            ub1=-4.1340125e-018            lub1=7.6318268e-025 wub1=-1.4293376e-024            pub1=1.5000638e-030             uc1=1.0453016e-009 luc1=-3.6705843e-016            wuc1=-1.6585434e-015            puc1=7.0669883e-022 at=70518.81                   lu0=2.06681e-010               pu0=8.1049318e-018 lpdiblc2=1.2689818e-009             wpdiblc2=3.8175403e-010             ppdiblc2=-3.4243337e-016 laigbinv=6.2548661e-011             paigbinv=1.8470289e-016             lbigc=-1.381539e-009 pbigc=1.5630361e-015             lbigsd=4.3547712e-010             pbigsd=-4.5387618e-016 lkt2=4.8042065e-009             pkt2=-4.2356854e-015            lute=6.5236608e-007 pute=-7.9661348e-013            lat=0.026444627                wat=0.044398672 pat=-3.9825608e-008            leta0=0                          weta0=0 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' ua1_ff=-9.96664e-11               ua1_ss=9.96664e-11                ua1_fs=9.96664e-11 ua1_sf=-9.96664e-11               lua1_ff=4.45512e-17                lua1_ss=-4.45512e-17 lua1_fs=-4.45512e-17               lua1_sf=4.45512e-17                wua1_ff=-2.6e-22 wua1_ss=2.6e-22                    wua1_fs=2.6e-22                    wua1_sf=-2.6e-22 pua1_ff=4.9e-28                    pua1_ss=-4.9e-28                   pua1_fs=-4.9e-28 pua1_sf=4.9e-28 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.3 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.46440048 lvth0=4.5305931e-009             wvth0=-3.7338203e-009            pvth0=1.2606295e-015 k2=0.028535487                lk2=-8.6307473e-010            wk2=-1.8656318e-008 pk2=-1.1817062e-015            cit=0.0049366722               lcit=-4.67281e-010 wcit=-3.372546e-009             pcit=6.2926306e-016             voff=-0.13781777 lvoff=-1.9708634e-010            wvoff=-9.2317988e-009            pvoff=3.5294159e-016 eta0=0.12                       etab=-0.05469247                wetab=-6.8228622e-008 u0=0.0096311878               wu0=7.6632907e-010             ua=3.017601e-010 lua=-3.6347071e-016            wua=-2.9869434e-016            pua=8.7419202e-023 ub=9.0351941e-019             lub=1.2357186e-025             wub=3.1773636e-025 pub=-1.0734814e-031            uc=3.7500961e-011             luc=-2.096473e-017 wuc=-1.9336799e-016            puc=2.5445201e-023             vsat=87550 wvsat=-0.0113703                 a0=2.398823                   la0=-3.3734649e-007 wa0=1.4715556e-007             pa0=-3.6259845e-014            ags=1.6792589 lags=-7.0345135e-008            wags=4.322408e-007              pags=-4.3629812e-014 keta=-0.072270513               lketa=-1.0294181e-008            wketa=6.1224692e-009 pketa=2.7758401e-014             pclm=-0.23865263                lpclm=1.8590003e-007 wpclm=2.972376e-007              ppclm=-9.8417893e-014            pdiblc2=0.0030377731 aigbacc=0.011475062                laigbacc=-2.414629e-011             waigbacc=2.3614192e-011 paigbacc=-1.9924055e-018            aigbinv=0.0073502416               waigbinv=3.1825824e-009 aigc=0.0044791455               laigc=3.8672285e-010             waigc=1.5671557e-009 paigc=-3.7231209e-016            bigc=-0.00035113353             wbigc=1.8482909e-009 aigsd=0.0053573032               laigsd=-7.371372e-011             waigsd=-4.3785235e-010 paigsd=1.1223663e-016             bigsd=0.00069325397              wbigsd=-5.1694048e-010 tvoff=0.000710187                ltvoff=3.38735e-010               wtvoff=1.47257e-009 ptvoff=-5.85184e-016              kt1=-0.2872798                 lkt1=1.5264275e-008 wkt1=9.040252e-008              pkt1=-2.7403017e-014            kt2=-0.086875474 wkt2=3.0707844e-008             ute=-0.90494786                wute=-2.9480272e-007 ua1=4.9007107e-009             lua1=-1.2054416e-015            wua1=-3.9602447e-015 pua1=1.0523549e-021             ub1=-6.6107367e-018            lub1=1.8702784e-024 wub1=5.4600511e-024             pub1=-1.5794929e-030            uc1=-1.181572e-010 luc1=1.5300763e-016             wuc1=1.4168702e-016             puc1=-9.8004151e-023 at=199558.92                  lu0=1.5532006e-010             pu0=-2.0633745e-016 lpdiblc2=-4.9777165e-010            wpdiblc2=-3.4319443e-009            ppdiblc2=1.3622898e-015 laigbinv=8.6738892e-010             paigbinv=-8.227181e-016             lbigc=4.3538986e-010 pbigc=-4.3412014e-016            lbigsd=-7.3113096e-011            pbigsd=1.1010832e-016 lkt2=1.1077621e-008             pkt2=-7.9602049e-015            lute=5.917323e-009 pute=6.4769602e-016             lat=-0.031236302               wat=-0.093400326 pat=2.1770544e-008             leta0=0                          weta0=0 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.4 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.44011074 lvth0=-6.4312113e-010            wvth0=-1.1916403e-009            pvth0=7.1914516e-016 k2=0.033498763                lk2=-1.9202526e-009            wk2=-3.138743e-008 pk2=1.5300207e-015             cit=0.0018134438               lcit=1.9796665e-010 wcit=-1.9239881e-010            pcit=-4.8108294e-017            voff=-0.11282517 lvoff=-5.5205096e-009            wvoff=-1.3319777e-008            pvoff=1.2236809e-015 eta0=0.12                       etab=-0.054692484               wetab=-6.822861e-008 u0=0.010497049                wu0=-3.4684829e-010            ua=-1.2577964e-009 lua=-3.1285163e-017            wua=1.1786562e-016             pua=-1.3080678e-024 ub=1.5309183e-018             lub=-1.0064104e-026            wub=-1.5798848e-025 pub=-6.0187488e-033            uc=-1.0010664e-010            luc=8.3456895e-018 wuc=-7.7506597e-017            puc=7.6672491e-025             vsat=87550 wvsat=-0.0113703                 a0=2.8317189                  la0=-4.2955331e-007 wa0=-1.577317e-007             pa0=2.868114e-014              ags=1.5899762 lags=-5.1327929e-008            wags=3.8442443e-007             pags=-3.3444925e-014 keta=0.00030238095              lketa=-2.5752207e-008            wketa=1.2074176e-007 pketa=3.3444925e-015             pclm=0.86924213                 lpclm=-5.0081549e-008 wpclm=-3.2819702e-007            ppclm=3.4799682e-014             pdiblc2=-0.0026198094 aigbacc=0.011121675                laigbacc=5.1125162e-011             waigbacc=7.0164038e-010 paigbacc=-1.4641198e-016            aigbinv=0.011021739                waigbinv=1.1978546e-010 aigc=0.0065854186               laigc=-6.1913297e-011            waigc=-5.8440546e-010 paigc=8.5970441e-017             bigc=0.002052715                wbigc=-7.0781466e-010 aigsd=0.0051419356               laigsd=-2.784042e-011             waigsd=-8.0699518e-011 paigsd=3.6163081e-017             bigsd=0.00060945333              wbigsd=-1.9784322e-010 tvoff=0.00305246                 ltvoff=-1.60169e-010              wtvoff=-1.93188e-009 ptvoff=1.39962e-016               kt1=-0.18801874                lkt1=-5.8783303e-009 wkt1=-5.3448551e-008            pkt1=3.2372607e-015             kt2=-0.0298104 wkt2=-1.5219152e-008            ute=-0.56660186                wute=-7.6030489e-007 ua1=-9.613096e-010             lua1=4.3168742e-017             wua1=1.1842544e-015 pua1=-4.3423382e-023            ub1=3.245131e-018              lub1=-2.2902139e-025 wub1=-2.9257673e-024            pub1=2.0668642e-031             uc1=9.7206034e-010 luc1=-7.9208704e-017            wuc1=-4.9433666e-016            puc1=3.7468893e-023 at=43763.095                  lu0=-2.9108377e-011            pu0=3.0769331e-017 lpdiblc2=7.0729341e-010             wpdiblc2=6.5803879e-009             ppdiblc2=-7.7033696e-016 laigbinv=8.5359995e-011             paigbinv=-1.7034236e-016            lbigc=-7.6629882e-011 pbigc=1.1033035e-016             lbigsd=-5.526356e-011             pbigsd=4.2140606e-017 lkt2=-1.0772401e-009            pkt2=1.8222452e-015             lute=-6.6150375e-008 pute=9.9799657e-014             lat=0.0019482085               wat=0.019400995 pat=-2.2561377e-009            letab=2.9531943e-015             petab=-2.675594e-021 leta0=0                          weta0=0                          peta0=0 lvsat=0                          pvsat=0                          jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)' jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                vsat_ff=4156.31 vsat_ss=-3465.84                   wvsat_ff=-0.00314005                wvsat_ss=0.00314005 lvsat_ff=-0.000885299               lvsat_ss=0.000738225                pvsat_ff=6.68834e-10 pvsat_ss=-6.68831e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.5 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.42788631 lvth0=-1.7066465e-009            wvth0=2.9273398e-009             pvth0=3.6079389e-016 k2=0.033586055                lk2=-1.927847e-009             wk2=-1.4013074e-008 pk2=1.8451708e-017             cit=0.0030041445               lcit=9.4375683e-011 wcit=-9.6103038e-010            pcit=1.8762652e-017             voff=-0.13225116 lvoff=-3.8304481e-009            wvoff=-7.1614406e-009            pvoff=6.8790566e-016 eta0=0.15799778                 etab=-0.069315496               wetab=-1.1021558e-007 u0=0.009669238                wu0=1.4319741e-009             ua=-1.7303953e-009 lua=9.8309403e-018             wua=2.5782619e-016             pua=-1.3484638e-023 ub=1.6606258e-018             lub=-2.1348653e-026            wub=-3.6584991e-025 pub=1.2065195e-032             uc=6.073366e-011              luc=-5.6474167e-018 wuc=-1.660097e-016             puc=8.4664945e-024             vsat=113952.62 wvsat=-0.037264888               a0=6.1133843                  la0=-7.150582e-007 wa0=-8.4564495e-007            pa0=8.8529593e-014             ags=1 lags=0                          wags=0                          pags=0 keta=0.43245916                 lketa=-6.3349847e-008            wketa=-3.46508e-007 pketa=4.3995221e-014             pclm=0.26740438                 lpclm=2.2783353e-009 wpclm=4.8045589e-008             ppclm=2.066575e-015              pdiblc2=0.0051629167 aigbacc=0.011516862                laigbacc=1.6743853e-011             waigbacc=-1.2376097e-009 paigbacc=2.2302777e-017             aigbinv=0.014877146                waigbinv=-4.4422508e-009 aigc=0.0068759793               laigc=-8.7192084e-011            waigc=-3.3064081e-010 paigc=6.3892917e-017             bigc=0.0022333419               wbigc=-3.1556754e-010 aigsd=0.0040626014               laigsd=6.6061656e-011             waigsd=8.6986872e-010 paigsd=-4.6536355e-017            bigsd=-0.00069235833             wbigsd=7.8265565e-010 tvoff=0.00226343                 ltvoff=-9.15232e-011              wtvoff=-2.66822e-009 ptvoff=2.04024e-016               kt1=-0.13640223                lkt1=-1.0368967e-008 wkt1=-2.2251562e-007            pkt1=1.7946096e-014             kt2=-0.045863333 wkt2=2.1556417e-008             ute=-1.2096085                 wute=2.805053e-007 ua1=-3.1058375e-009            lua1=2.2974267e-016             wua1=5.3457885e-015 pua1=-4.0547685e-022            ub1=4.3502045e-018             lub1=-3.2516279e-025 wub1=-6.8508875e-024            pub1=5.4817188e-031             uc1=5.4461334e-010 luc1=-4.2020815e-017            wuc1=-7.8794907e-016            puc1=6.3013173e-023 at=62469.172                  lu0=4.2911183e-011             pu0=-1.2398821e-016 lpdiblc2=3.019625e-011              wpdiblc2=-3.8848525e-009            ppdiblc2=1.4013895e-016 laigbinv=-2.5006047e-010            paigbinv=2.2655479e-016             lbigc=-9.2344419e-011 pbigc=7.6204855e-017             lbigsd=5.7994055e-011             pbigsd=-4.3162796e-017 lkt2=3.1936514e-010             pkt2=-1.3772293e-015            lute=-1.0208797e-008 pute=9.2491705e-015             lat=0.00032077988              wat=0.035160335 pat=-3.6272003e-009            letab=1.272205e-009              petab=3.652864e-015 leta0=-3.3058069e-009            weta0=4.8433921e-010             peta0=-4.2137511e-017 lvsat=-0.0022970275              pvsat=2.2528292e-009 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=-13841.5                   vsat_ss=12130.4                    wvsat_ff=0.0116345 wvsat_ss=-0.0109902                 ua1_ff=1.06941e-10                lua1_ff=-9.30382e-18 wua1_ff=-1.61063e-16               pua1_ff=1.40125e-23                lvsat_ff=0.000680518 lvsat_ss=-0.000618653               pvsat_ff=-6.16549e-10               pvsat_ss=5.605e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.6 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.41326458 lvth0=-2.4523546e-009            wvth0=-1.1864992e-008            pvth0=1.1152029e-015 k2=0.11518119                 lk2=-6.0891986e-009            wk2=-6.1047269e-008 pk2=2.4171956e-015             cit=0.0071767386               lcit=-1.1842662e-010 wcit=-4.5777092e-009            pcit=2.0321327e-016             voff=-0.12383233 lvoff=-4.2598086e-009            wvoff=-2.6072682e-008            pvoff=1.652379e-015 eta0=0.003466172                etab=0.066954387                wetab=-1.6889898e-007 u0=0.0089749473               wu0=1.4955035e-009             ua=-3.1298798e-009 lua=8.1204647e-017             wua=1.1902163e-015             pua=-6.1036534e-023 ub=3.6189063e-018             lub=-1.2122096e-025            wub=-1.9553395e-024 pub=9.3129163e-032             uc=3.7736097e-010             luc=-2.1795409e-017 wuc=-3.8718904e-016            puc=1.9746641e-023             vsat=34969.068 wvsat=0.043401609                a0=0.5730515                  la0=-4.3250123e-007 wa0=1.1548367e-005             pa0=-5.4356502e-013            ags=1 lags=0                          wags=0                          pags=0 keta=-2.2750033                 lketa=7.4730739e-008             wketa=2.181953e-006 pketa=-8.4956289e-014            pclm=0.20007811                 lpclm=5.7119751e-009 wpclm=1.6644017e-007             ppclm=-3.9715488e-015            pdiblc2=0.0046116667 aigbacc=0.014086504                laigbacc=-1.1430786e-010            waigbacc=-4.0956903e-009 paigbacc=1.6806489e-016             aigbinv=0.009974                   aigc=0.0030539549 laigc=1.0773116e-010             waigc=3.808172e-009              paigc=-1.4718654e-016 bigc=-0.0026760174              wbigc=5.0561602e-009             aigsd=0.0064797994 laigsd=-5.7215443e-011            waigsd=-1.054352e-009             paigsd=5.1598901e-017 bigsd=0.0017646767               wbigsd=-1.2151061e-009            tvoff=-0.00197831 ltvoff=1.24805e-010               wtvoff=2.45895e-009               ptvoff=-5.74619e-017 kt1=-0.52020817                lkt1=9.2051363e-009             wkt1=1.4538834e-007 pkt1=-8.1700597e-016            kt2=-0.10257763                wkt2=2.4322891e-008 ute=2.5720197                  wute=-4.8368498e-006            ua1=1.060051e-008 lua1=-4.6928106e-016            wua1=-9.8990411e-015            pua1=3.7200946e-022 ub1=-1.1193374e-017            lub1=4.6755969e-025             wub1=1.0412782e-023 pub1=-3.3227529e-031            uc1=1.0658057e-009             luc1=-6.8601627e-017 wuc1=5.9144847e-017             puc1=1.9811383e-023             at=174212.15 lu0=7.8320011e-011             pu0=-1.2722821e-016            lpdiblc2=5.831e-011 wpdiblc2=-6.44317e-009              ppdiblc2=2.7061314e-016             lbigc=1.580329e-010 pbigc=-1.9775326e-016            lbigsd=-6.731473e-011             pbigsd=5.8723051e-017 lkt2=3.2117944e-009             pkt2=-1.5183195e-015            lute=-2.0307183e-007 pute=2.7023428e-013             lat=-0.0053781118              wat=-0.13060577 pat=4.8268712e-009             letab=-5.677559e-009             petab=6.6457175e-015 leta0=4.5753051e-009             weta0=6.268226e-008              peta0=-3.2142315e-015 lvsat=0.0017311334               pvsat=-1.8611622e-009 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=-2822.26                   wvsat_ff=-0.00257705                ua1_ff=-4.27762e-10 ua1_ss=-1.4091e-10                lua1_ff=1.7966e-17                 lua1_ss=7.1864e-18 wua1_ff=6.44252e-16                wua1_ss=2.12224e-16                pua1_ff=-2.70586e-23 pua1_ss=-1.08234e-23               lvsat_ff=0.000118536                pvsat_ff=1.08234e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.7 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.47315579 lvth0=6.307568e-011              wvth0=5.2307089e-009             pvth0=3.9718333e-016 k2=0.10984405                 lk2=-5.865039e-009             wk2=-5.1022422e-008 pk2=1.9961521e-015             cit=-0.008586102               lcit=5.4361269e-010 wcit=4.7691274e-009             pcit=-1.8935387e-016            voff=-0.23863808 lvoff=5.6203289e-010             wvoff=5.2783865e-008             pvoff=-1.659596e-015 eta0=0.0018443259               etab=-0.14252098                wetab=-7.7078619e-008 u0=0.024229534                wu0=-1.3753818e-008            ua=-4.1929381e-010 lua=-3.2639964e-017            wua=-2.1094213e-015            pua=7.7548244e-023 ub=5.8554529e-019             lub=6.1802032e-027             wub=1.8649834e-024 pub=-6.7324397e-032            uc=4.803526e-011              luc=-7.9637296e-018 wuc=-7.7983582e-017            puc=6.7600118e-024             vsat=60305.67 wvsat=-0.0010682456              a0=11.763408                  la0=-9.0249621e-007 wa0=-1.0464818e-005            pa0=3.8098877e-013             ags=1 lags=0                          wags=0                          pags=0 keta=-0.30895667                lketa=-7.84322e-009              wketa=6.3446274e-007 pketa=-1.9961699e-014            pclm=0.51258252                 lpclm=-7.4132101e-009 wpclm=5.7911303e-009             ppclm=2.775711e-015              pdiblc2=0.0023333333 aigbacc=0.0075896422               laigbacc=1.5856033e-010             waigbacc=5.8370631e-009 paigbacc=-2.4911076e-016            aigbinv=0.009974                   aigc=0.0058257731 laigc=-8.6852034e-012            waigc=6.6650185e-010             paigc=-1.523639e-017 bigc=0.00095663003              wbigc=1.1636008e-009             aigsd=0.0047004023 laigsd=1.7519234e-011             waigsd=3.6576287e-010             paigsd=-8.0459234e-018 bigsd=-0.00010965818             wbigsd=2.2488322e-010             tvoff=0.00343845 ltvoff=-1.02699e-010              wtvoff=3.73405e-010               ptvoff=3.01311e-017 kt1=-0.40321064                lkt1=4.2912397e-009             wkt1=3.7520552e-007 pkt1=-1.0469328e-014            kt2=-0.0021925248              wkt2=-4.7507191e-008 ute=-8.7274453                 wute=7.4540655e-006             ua1=6.9177738e-009 lua1=-3.1460613e-016            wua1=-7.072747e-015             pua1=2.5330511e-022 ub1=-1.4794301e-017            lub1=6.1879865e-025             wub1=1.3818018e-023 pub1=-4.7529517e-031            uc1=-1.8304025e-009            luc1=5.3039119e-017 wuc1=1.599174e-015              puc1=-4.486984e-023             at=-29400.689 lu0=-5.6237266e-010            pu0=5.1324328e-016             lpdiblc2=1.54e-010 lbigc=5.4617121e-012             pbigc=-3.4265765e-017            lbigsd=1.1407333e-011 pbigsd=-1.7564982e-018            lkt2=-1.0043801e-009            pkt2=1.4985439e-015 lute=2.715057e-007              pute=-2.4598416e-013            lat=0.0031736273 wat=0.035289252                pat=-2.1407199e-009            letab=3.1204063e-009 petab=2.7892622e-015             leta0=4.6434227e-009             weta0=-3.094173e-008 peta0=7.1797611e-016             lvsat=0.00066699613              pvsat=6.5717064e-012 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' voff_ff=0.0110715                  voff_ss=-0.0166072                 voff_mcl=-0.0256667 lvoff_ff=-4.65003e-10               lvoff_ss=6.97504e-10                lvoff_mcl=1.078e-09 wvoff_ff=-1.66748e-08               wvoff_ss=2.50122e-08                wvoff_mcl=1.1e-14 pvoff_ff=7.0034e-16                 pvoff_ss=-1.05051e-15               pvoff_mcl=9e-22 u0_ff=-0.000276787               u0_ss=0.000276787                wu0_ff=4.16869e-10 wu0_ss=-4.16869e-10               vsat_ff=-2767.87                   vsat_sf=-8267.86 vsat_fs=7333.31                    wvsat_ff=0.00416869                 wvsat_sf=0.00416872 wvsat_fs=-3.2e-08                   ua1_ss=1.4091e-10                 lua1_ss=-4.65003e-18 wua1_ss=-2.12224e-16               pua1_ss=7.0034e-24                 lu0_ff=1.16251e-11 lu0_ss=-1.16251e-11               pu0_ff=-1.75085e-17               pu0_ss=1.75085e-17 lvsat_ff=0.000116251                lvsat_sf=0.000347251                lvsat_fs=-0.000308001 pvsat_ff=-1.75085e-10               pvsat_sf=-1.75085e-10               pvsat_fs=-2.6e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_hvt_mac.8 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.50792064 lvth0=3.3491036e-008             wvth0=1.1793879e-008             pvth0=-7.1886426e-015 k2=0.020092527                lk2=3.0042411e-009             wk2=-1.5543174e-008 pk2=2.6571405e-015             cit=0.0015972017               lcit=-6.0518517e-014 wcit=-2.015829e-010             pcit=2.1863939e-020             voff=-0.14599861 lvoff=-2.0563679e-012            wvoff=-5.0839813e-010            pvoff=-1.6976383e-019 eta0=0.12                       etab=-0.067043167               wetab=-5.7038891e-008 u0=0.010003233                wu0=6.32086e-011               ua=-2.8237273e-010 lua=-1.7435648e-016            wua=1.6580668e-016             pua=-1.6158398e-023 ub=1.6107658e-018             lub=1.9457319e-026             wub=-3.0018046e-025 pub=1.1830486e-033             uc=-5.5052362e-010            luc=4.5456098e-016 wuc=1.1260495e-017             puc=-1.0131067e-022            vsat=52250 wvsat=0.0206115                  a0=1.5474191                  la0=4.0761703e-012 wa0=1.4885658e-007             pa0=-2.9708671e-018            ags=1.0047006 lags=6.0819066e-007             wags=-1.3325985e-007            pags=-8.5688772e-014 keta=-0.53851388                lketa=3.1801888e-007             wketa=1.8497281e-007 pketa=-5.7039278e-014            pclm=0.092778391                lpclm=-1.1015474e-011 wpclm=3.774565e-008              ppclm=7.8858038e-018             pdiblc2=0.0005 aigbacc=0.011745844                laigbacc=-1.1761774e-010            waigbacc=2.5897778e-010 paigbacc=3.4759966e-017             aigbinv=0.00986785                 waigbinv=5.482659e-010 aigc=0.0053537192               laigc=4.9830268e-011             waigc=3.8806773e-010 paigc=-2.1477384e-017            bigc=0.00072997667              wbigc=4.3064294e-010 aigsd=0.0052173076               laigsd=9.8022703e-016             waigsd=-1.4857026e-010 paigsd=9.5834417e-023             bigsd=0.00051797083              wbigsd=-1.9340457e-010 tvoff=0.0035215                  ltvoff=-2.17246e-009              wtvoff=-5.83141e-010 ptvoff=7.7119e-016                kt1=-0.16236379                lkt1=-7.5571552e-008 wkt1=-1.7291372e-008            pkt1=3.0782614e-014             kt2=-0.017666667 wkt2=-2.7482e-008               ute=-0.56826083                wute=-3.5568579e-007 ua1=3.616927e-009              lua1=2.3276875e-016             wua1=-8.832024e-016 pua1=-1.2709275e-022            ub1=-3.0976823e-018            lub1=-1.1059312e-029 wub1=7.4901278e-026             pub1=8.214379e-036              uc1=2.2250296e-009 luc1=-2.740378e-015             wuc1=-4.8031989e-016            puc1=8.4131614e-022 at=100000                     lu0=0                          pu0=0 lat=0                          wat=0                          pat=0 leta0=0                          weta0=0                          peta0=0 lvsat=0                          pvsat=0                          jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)' jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                ua1_ff=5.53022e-12 ua1_ss=-5.53022e-12               ua1_fs=-5.53022e-12               ua1_sf=5.53022e-12 lua1_ff=-4.98109e-17               lua1_ss=4.98109e-17                lua1_fs=4.98109e-17 lua1_sf=-4.98109e-17               wua1_ff=1e-24                      wua1_ss=-1e-24 wua1_fs=-1e-24                     wua1_sf=1e-24                      pua1_ff=-4.3e-29 pua1_ss=4.3e-29                    pua1_fs=4.3e-29                    pua1_sf=-4.3e-29 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.9 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.4905315 lvth0=1.7892971e-008             wvth0=1.1827956e-008             pvth0=-7.2192094e-015 k2=0.034008292                lk2=-9.4782001e-009            wk2=-1.6339827e-008 pk2=3.371738e-015              cit=0.00092279805              lcit=6.0487958e-010 wcit=9.6217185e-011             pcit=-2.6710481e-016            voff=-0.14695084 lvoff=8.5209699e-010             wvoff=1.2651117e-009             pvoff=-1.5910081e-015 eta0=0.12                       etab=-0.067043167               wetab=-5.7038891e-008 u0=0.0097809253               wu0=4.6829328e-011             ua=-2.6405512e-010 lua=-1.9078737e-016            wua=2.3549663e-016             pua=-7.8670282e-023 ub=1.8882463e-018             lub=-2.2944271e-025            wub=-4.973186e-025 pub=1.7801596e-031             uc=-1.8701556e-011            luc=-2.2483405e-017 wuc=-1.2079255e-016            puc=1.7140908e-023             vsat=52250 wvsat=0.0206115                  a0=0.93885832                 la0=5.4588305e-007 wa0=6.9544272e-007             pa0=-4.9029074e-013            ags=0.42968418 lags=1.1239804e-006             wags=4.9155339e-007             pags=-6.4614625e-013 keta=-0.26950075                lketa=7.6714104e-008             wketa=1.7186888e-007 pketa=-4.5285055e-014            pclm=-0.048211683               lpclm=1.2645708e-007 wpclm=5.0418349e-008             ppclm=-1.1359525e-014            pdiblc2=-6.3400042e-005 aigbacc=0.011816054                laigbacc=-1.8059616e-010            waigbacc=5.6633773e-010 paigbacc=-2.4094191e-016            aigbinv=0.0077674963               waigbinv=2.1820983e-009 aigc=0.0041783814               laigc=1.1041083e-009             waigc=1.1701333e-009 paigc=-7.2299016e-016            bigc=-0.00070638499             wbigc=1.384872e-009 aigsd=0.0056410187               laigsd=-3.8006787e-010            waigsd=-4.7209162e-010 paigsd=2.9019876e-016             bigsd=0.00098230864              wbigsd=-5.4794757e-010 tvoff=0.000268003                ltvoff=7.45926e-010               wtvoff=8.10886e-010 ptvoff=-4.79252e-016              kt1=-0.29307346                lkt1=4.1675022e-008 wkt1=5.2993676e-008             pkt1=-3.2263074e-014            kt2=-0.0011084614 wkt2=-4.2614086e-008            ute=0.27774709                 wute=-8.9299415e-007 ua1=9.9029022e-009             lua1=-5.405751e-015             wua1=-4.4025192e-015 pua1=3.0297344e-021             ub1=-9.3457973e-018            lub1=5.6045481e-024 wub1=3.2925395e-024             pub1=-2.8862132e-030            uc1=-2.1788866e-009 luc1=1.2099349e-015             wuc1=1.2625711e-015             puc1=-7.2205711e-022 at=149135.32                  lu0=1.9941028e-010             pu0=1.4692207e-017 lpdiblc2=5.0536984e-010             wpdiblc2=-3.8951956e-010            ppdiblc2=3.4939905e-016 laigbinv=1.8840172e-009             paigbinv=-1.4655477e-015            lbigc=1.2884164e-009 pbigc=-8.5594349e-016            lbigsd=-4.1651101e-010            pbigsd=3.1802506e-016 lkt2=-1.485271e-008             pkt2=1.3573481e-014             lute=-7.5886911e-007 pute=4.8196561e-013             lat=-0.044074379               wat=-0.026827883 pat=2.4064611e-008             leta0=0                          weta0=0 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' ua1_ff=-9.96669e-11               ua1_ss=9.96669e-11                ua1_fs=9.96669e-11 ua1_sf=-1.74995e-10               lua1_ff=4.4551e-17                 lua1_ss=-4.4551e-17 lua1_fs=-4.4551e-17                lua1_sf=1.1212e-16                 wua1_ff=3e-23 wua1_ss=-3e-23                     wua1_fs=-3e-23                     wua1_sf=6.8247e-17 pua1_ff=2.9e-29                    pua1_ss=-2.9e-29                   pua1_fs=-2.9e-29 pua1_sf=-6.12175e-23 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.10 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.46045486 lvth0=4.4487166e-009             wvth0=-7.3085519e-009            pvth0=1.3348097e-015 k2=0.018452575                lk2=-2.5247942e-009            wk2=-9.5211998e-009 pk2=3.2381163e-016             cit=0.0019688546               lcit=1.3729232e-010 wcit=-6.8370328e-010            pcit=8.1519636e-017             voff=-0.14912272 lvoff=1.8229284e-009             wvoff=1.0104892e-009             pvoff=-1.4771918e-015 eta0=0.12                       etab=-0.067043167               wetab=-5.7038891e-008 u0=0.010719012                wu0=-2.1923942e-010            ua=-1.3933474e-010 lua=-2.4653738e-016            wua=1.0093759e-016             pua=-1.8522392e-023 ub=1.5087024e-018             lub=-5.9786592e-026            wub=-2.3055946e-025 pub=5.877462e-032              uc=-5.3866987e-011            luc=-6.7644567e-018 wuc=-1.1058862e-016            puc=1.2579753e-023             vsat=52250 wvsat=0.0206115                  a0=3.6628141                  la0=-6.7172518e-007 wa0=-9.9802034e-007            pa0=2.6668725e-013             ags=2.7431297 lags=8.9870288e-008             wags=-5.3162616e-007            pags=-1.8878499e-013 keta=-0.21428518                lketa=5.2032744e-008             wketa=1.3478776e-007 pketa=-2.8709793e-014            pclm=0.16462378                 lpclm=3.1319627e-008 wpclm=-6.8130824e-008            ppclm=4.1631956e-014             pdiblc2=-0.0030710769 aigbacc=0.011463599                laigbacc=-2.304882e-011             waigbacc=3.399948e-011 paigbacc=-2.986713e-018             aigbinv=0.011109836                waigbinv=-2.2361011e-010 aigc=0.0072027777               laigc=-2.4779691e-010            waigc=-9.0045506e-010 paigc=2.0256282e-016             bigc=0.002859286                wbigc=-1.0603492e-009 aigsd=0.004326946                laigsd=2.0732264e-010             waigsd=4.9565126e-010 paigsd=-1.4238231e-016            bigsd=-0.00047818301             wbigsd=5.4438143e-010 tvoff=0.00306691                 ltvoff=-5.05185e-010              wtvoff=-6.62625e-010 ptvoff=1.79407e-016               kt1=-0.14700798                lkt1=-2.3616247e-008 wkt1=-3.668375e-008             pkt1=7.8227353e-015             kt2=-0.031573792 wkt2=-1.939548e-008             ute=-1.5380494                 wute=2.7878727e-007 ua1=-3.3793506e-009            lua1=5.3141598e-016             wua1=3.5414908e-015 pua1=-5.2123803e-022            ub1=4.3341616e-018             lub1=-5.1039351e-025 wub1=-4.4560268e-024            pub1=5.7739587e-031             uc1=3.5186139e-010 luc1=7.8690513e-017             wuc1=-2.8414982e-016            puc1=-3.0672841e-023 at=91111.267                  lu0=-2.1991435e-010            pu0=1.3362494e-016 lpdiblc2=1.8498014e-009             wpdiblc2=2.1026738e-009             ppdiblc2=-7.6461139e-016 laigbinv=3.8999144e-010             paigbinv=-3.9019599e-016            lbigc=-3.0543852e-010 pbigc=2.3707038e-016             lbigsd=2.3632876e-010             pbigsd=-1.70246e-016 lkt2=-1.2347073e-009            pkt2=3.1947643e-015             lute=5.2791923e-008 pute=-4.1820691e-014            lat=-0.018137629               wat=0.0048532481 pat=9.9031453e-009             leta0=0                          weta0=0 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' ua1_sf=1.44861e-10                lua1_sf=-3.08554e-17               wua1_sf=-1.31244e-16 pua1_sf=2.7955e-23 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.11 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.43272224 lvth0=-1.4583313e-009            wvth0=-7.8856218e-009            pvth0=1.4577256e-015 k2=0.0090062369               lk2=-5.1272428e-010            wk2=-9.1972018e-009 pk2=2.5480007e-016             cit=0.0018964851               lcit=1.5270701e-010 wcit=-2.6763429e-010            pcit=-7.1030589e-018            voff=-0.11562867 lvoff=-5.311305e-009             wvoff=-1.0779808e-008            pvoff=1.0341415e-015 eta0=0.12                       etab=-0.067043167               wetab=-5.7038891e-008 u0=0.0091998449               wu0=8.2841872e-010             ua=-1.2119961e-009 lua=-1.8060505e-017            wua=7.6370528e-017             pua=-1.3289608e-023 ub=1.3096514e-018             lub=-1.7388713e-026            wub=4.2479385e-026 pub=6.1734713e-034             uc=-8.4073845e-011            luc=-3.3039596e-019 wuc=-9.203231e-017             puc=8.6272584e-024             vsat=52250 wvsat=0.0206115                  a0=2.3689586                  la0=-3.9613396e-007 wa0=2.6152916e-007             pa0=-1.596793e-015             ags=4.6599755 lags=-3.1841787e-007            wags=-2.3969949e-006            pags=2.0853856e-013 keta=0.21364937                 lketa=-3.9117316e-008            wketa=-7.2550615e-008 pketa=1.5453281e-014             pclm=0.26401306                 lpclm=1.014971e-008 wpclm=2.2014051e-007             ppclm=-1.9769839e-014            pdiblc2=0.0074179525 aigbacc=0.011734578                laigbacc=-8.0767214e-011            waigbacc=1.4635055e-010 paigbacc=-2.6917491e-017            aigbinv=0.014989274                waigbinv=-3.4748012e-009 aigc=0.0056407277               laigc=8.4919748e-011             waigc=2.7148445e-010 paigc=-4.7060298e-017            bigc=0.00089707029              wbigc=3.3919947e-010 aigsd=0.0053767296               laigsd=-1.6281262e-011            waigsd=-2.9342289e-010 paigsd=2.5690484e-017             bigsd=0.00085935417              wbigsd=-4.2425338e-010 tvoff=0.000490776                ltvoff=4.35316e-011               wtvoff=3.89007e-010 ptvoff=-4.45906e-017              kt1=-0.24587845                lkt1=-2.556836e-009 wkt1=-1.0276543e-009            pkt1=2.2798697e-016             kt2=-0.049603245 wkt2=2.7131661e-009             ute=-1.7300069                 wute=2.9374005e-007 ua1=-1.4715999e-009            lua1=1.250651e-016              wua1=1.6465774e-015 pua1=-1.1762148e-022            ub1=2.6313832e-018             lub1=-1.477017e-025 wub1=-2.3697118e-024            pub1=1.3301078e-031             uc1=1.2234099e-009 luc1=-1.0694932e-016            wuc1=-7.2205934e-016            puc1=6.2601886e-023 at=-20025.154                 lu0=1.036682e-010              pu0=-8.9526247e-017 lpdiblc2=-3.8436186e-010            wpdiblc2=-2.5138243e-009            ppdiblc2=2.1870272e-016 laigbinv=-4.3632882e-010            paigbinv=3.023077e-016              lbigc=1.1251342e-010 pbigc=-6.103348e-017             lbigsd=-4.8566663e-011            pbigsd=3.6073217e-017 lkt2=2.6055663e-009             pkt2=-1.5143773e-015            lute=9.3678862e-008 pute=-4.5005632e-014            lat=0.0055344289               wat=0.077193148 pat=-5.5052534e-009            leta0=0                          weta0=0 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=690.478                    wvsat_ff=3.3e-10                    ua1_fs=5.23611e-11 lua1_fs=-1.11529e-17               wua1_fs=-4.74392e-17               pua1_fs=1.01045e-23 lvsat_ff=-0.000147072               pvsat_ff=1.5e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.12 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.4253388 lvth0=-2.1006905e-009            wvth0=6.1929565e-010             pvth0=7.1779774e-016 k2=0.016326971                lk2=-1.1496282e-009            wk2=1.6236556e-009 pk2=-6.8661453e-016            cit=0.0015575356               lcit=1.8219562e-010 wcit=3.4959731e-010             pcit=-6.0802208e-017            voff=-0.12961119 lvoff=-4.0948251e-009            wvoff=-9.553253e-009             pvoff=9.2743122e-016 eta0=0.1877569                  etab=-0.13128605                wetab=-5.4070263e-008 u0=0.01239785                 wu0=-1.0401487e-009            ua=-8.4795558e-010 lua=-4.9732033e-017            wua=-5.4166423e-016            pua=4.0479416e-023 ub=5.6600755e-019             lub=4.7308298e-026             wub=6.258742e-025 pub=-5.0138002e-032            uc=-2.4987725e-010            luc=1.40945e-017 wuc=1.1540379e-016             puc=-9.4196822e-024            vsat=25605.075 wvsat=0.042777983                a0=6.9226118                  la0=-7.9230179e-007 wa0=-1.578805e-006             pa0=1.5851228e-013             ags=1 lags=0                          wags=0                          pags=0 keta=0.32621748                 lketa=-4.8910742e-008            wketa=-2.5025304e-007 pketa=3.0913392e-014             pclm=0.27674632                 lpclm=9.0419167e-009 wpclm=3.9581785e-008             ppclm=-4.0612298e-015            pdiblc2=0.000875 aigbacc=0.009990163                laigbacc=7.0996859e-011             waigbacc=1.4557993e-010 paigbacc=-2.6850447e-017            aigbinv=0.009974                   aigc=0.0065427893 laigc=6.4403892e-012             waigc=-2.8770652e-011            paigc=-2.0938104e-017 bigc=0.0019213177               wbigc=-3.287364e-011             aigsd=0.0049059217 laigsd=2.4679022e-011             waigsd=1.0582048e-010             paigsd=-9.0436892e-018 bigsd=5.2531917e-005             wbigsd=1.0778508e-010             tvoff=-0.00207596 ltvoff=2.66838e-010               wtvoff=1.26327e-009               ptvoff=-1.20651e-016 kt1=-0.51401059                lkt1=2.077066e-008              wkt1=1.1959755e-007 pkt1=-1.0266406e-014            kt2=-0.0021444762              wkt2=-1.8052867e-008 ute=-0.58405306                wute=-2.8624793e-007            ua1=4.8571094e-009 lua1=-4.2553261e-016            wua1=-1.8686414e-015            pua1=1.8820256e-022 ub1=-5.3745143e-018            lub1=5.4881138e-025             wub1=1.9597078e-024 pub1=-2.4364873e-031            uc1=-5.2997649e-010            luc1=4.5595299e-017 wuc1=1.8562932e-016             puc1=-1.6367027e-023            at=109042.77 lu0=-1.7455828e-010            pu0=7.3039119e-017             lpdiblc2=1.84875e-010 lbigc=2.3403897e-011             pbigc=-2.8663119e-017            lbigsd=2.1626873e-011 pbigsd=-1.0214129e-017            lkt2=-1.5233466e-009            pkt2=2.9226752e-016 lute=-6.0191192e-009            pute=5.453322e-015              lat=-0.0056944803 wat=-0.0070353442              pat=1.8226254e-009             letab=5.5891307e-009 petab=-2.5827068e-016            leta0=-5.89485e-009              weta0=-2.647742e-008 peta0=2.3035355e-015             lvsat=0.0023181084               pvsat=-1.928484e-009 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=1148.62                    wvsat_ff=-0.00194664                ua1_ff=-1.78264e-10 ua1_ss=1.07431e-10                ua1_fs=-7.58334e-11               lua1_ff=1.5509e-17 lua1_ss=-9.34646e-18               lua1_fs=1.7e-24                    wua1_ff=9.73321e-17 wua1_ss=-9.73321e-17               wua1_fs=6.87049e-17                pua1_ff=-8.46789e-24 pua1_ss=8.46789e-24                pua1_fs=1.3e-30                    lvsat_ff=-0.000186929 pvsat_ff=1.69358e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.13 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.42156554 lvth0=-2.2931269e-009            wvth0=-4.344327e-009             pvth0=9.709425e-016 k2=0.085036785                lk2=-4.6538287e-009            wk2=-3.3736442e-008 pk2=1.1167505e-015             cit=0.0060412492               lcit=-4.6473777e-011 wcit=-3.5489558e-009            pcit=1.38024e-016               voff=-0.14881809 lvoff=-3.1152737e-009            wvoff=-3.4355889e-009            pvoff=6.1543036e-016 eta0=-0.058930954               etab=0.11920697                 wetab=-2.1623983e-007 u0=0.0066518622               wu0=3.6002185e-009             ua=-2.4789848e-009 lua=3.3450455e-017             wua=6.0050543e-016             pua=-1.7771237e-023 ub=1.866857e-018              lub=-1.9035023e-026            wub=-3.6798282e-025 pub=5.4870622e-034             uc=1.710845e-010              luc=-7.374549e-018 wuc=-2.0030256e-016            puc=6.6813414e-024             vsat=60094.374 wvsat=0.02063808                 a0=11.868268                  la0=-1.0445302e-006 wa0=1.3149013e-006             pa0=1.0933258e-014             ags=1 lags=0                          wags=0                          pags=0 keta=-0.33733889                lketa=-1.5069367e-008            wketa=4.2642903e-007 pketa=-3.5973938e-015            pclm=0.8109853                  lpclm=-1.8204271e-008 wpclm=-3.8704174e-007            ppclm=1.769657e-014              pdiblc2=-0.016655556 aigbacc=0.015696705                laigbacc=-2.2003679e-010            waigbacc=-5.5545327e-009 paigbacc=2.638553e-016              aigbinv=0.009974                   aigc=0.008275614 laigc=-8.1933669e-011            waigc=-9.2265113e-010            paigc=2.46498e-017 bigc=0.0044923244               wbigc=-1.4383575e-009            aigsd=0.0062423777 laigsd=-4.3480235e-011            waigsd=-8.3924799e-010            paigsd=3.9154803e-017 bigsd=0.00090291122              wbigsd=-4.3434657e-010            tvoff=0.00492004 ltvoff=-8.99585e-011              wtvoff=-3.79095e-009              ptvoff=1.37114e-016 kt1=-0.053317342               lkt1=-2.7246956e-009            wkt1=-2.7761476e-007 pkt1=9.9914218e-015             kt2=-0.10404634                wkt2=2.5653543e-008 ute=-1.6450917                 wute=-1.016147e-006             ua1=-7.9588925e-009 lua1=2.2808348e-016             wua1=6.9157777e-015             pua1=-2.5980281e-022 ub1=1.3676794e-017             lub1=-4.2280536e-025            wub1=-1.211959e-023 pub1=4.7439545e-031             uc1=2.4082156e-009             luc1=-1.042525e-016 wuc1=-1.1570784e-015            puc1=5.2111069e-023             at=-124342.1 lu0=1.1848711e-010             pu0=-1.6361961e-016            lpdiblc2=1.0789333e-009 wpdiblc2=1.2824933e-008             ppdiblc2=-6.540716e-016             lbigc=-1.0771745e-010 pbigc=4.3016559e-017             lbigsd=-2.1742471e-011            pbigsd=1.7434585e-017 lkt2=3.6736485e-009             pkt2=-1.9367594e-015            lute=4.809385e-008 pute=4.2678172e-014             lat=0.0062081479               wat=0.13988437 pat=-5.6702801e-009            letab=-7.1860133e-009            petab=8.0123771e-015 leta0=6.6862304e-009             weta0=1.1921406e-007             peta0=-5.1267298e-015 lvsat=0.00055915418              pvsat=-7.9934898e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=-7183.32                   vsat_ss=-7077.78                   wvsat_ff=0.0013741 wvsat_ss=0.00641247                 ua1_ff=7.13056e-10                ua1_ss=-1.94833e-10 ua1_fs=-4.29722e-10               lua1_ff=-2.99483e-17               lua1_ss=6.06903e-18 lua1_fs=1.80483e-17                wua1_ff=-3.89328e-16               wua1_ss=2.61079e-16 wua1_fs=3.89328e-16                pua1_ff=1.63518e-23                pua1_ss=-9.81107e-24 pua1_fs=-1.63518e-23               lvsat_ff=0.000238                   lvsat_ss=0.000360967 pvsat_ff=-2e-16                     pvsat_ss=-3.27036e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.14 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.53228605 lvth0=2.3571345e-009             wvth0=5.8802731e-008             pvth0=-1.681234e-015 k2=0.10745595                 lk2=-5.5954337e-009            wk2=-4.8858805e-008 pk2=1.7518897e-015             cit=-0.0068143528              lcit=4.9346151e-010 wcit=3.1639227e-009             pcit=-1.439169e-016             voff=-0.22196328 lvoff=-4.317544e-011             wvoff=3.7676497e-008             pvoff=-1.1112773e-015 eta0=-0.020870132               etab=-0.089575945               wetab=-1.2504682e-007 u0=0.0044866296               wu0=4.133254e-009              ua=-4.6772524e-009 lua=1.257777e-016              wua=1.7482893e-015             pua=-6.5978158e-023 ub=5.2124826e-018             lub=-1.595513e-025             wub=-2.3270218e-024 pub=8.2828343e-032             uc=1.6471221e-010             luc=-7.1069126e-018 wuc=-1.8369289e-016            puc=5.9837356e-024             vsat=77334.321 wvsat=-0.016496204               a0=5.4045516                  la0=-7.7305416e-007 wa0=-4.7036943e-006            pa0=2.6371427e-013             ags=1 lags=0                          wags=0                          pags=0 keta=-0.64101111                lketa=-2.3151333e-009            wketa=9.3530407e-007 pketa=-2.4970145e-014            pclm=0.69167227                 lpclm=-1.3193124e-008 wpclm=-1.5646418e-007            ppclm=8.0123125e-015             pdiblc2=-0.002975 aigbacc=0.011061059                laigbacc=-2.5339645e-011            waigbacc=2.6919596e-009 paigbacc=-8.2497381e-017            aigbinv=0.016074539                waigbinv=-5.5270882e-009 aigc=0.0087925403               laigc=-1.0364457e-010            waigc=-2.0213892e-009 paigc=7.0796799e-017             bigc=0.0048280578               wbigc=-2.3439127e-009 aigsd=0.0036666661               laigsd=6.4699653e-011             waigsd=1.3023279e-009 paigsd=-5.0791383e-017            bigsd=-0.00076604748             wbigsd=8.1957193e-010 tvoff=0.00786928                 ltvoff=-2.13826e-010              wtvoff=-3.64092e-009 ptvoff=1.30813e-016               kt1=0.44304802                 lkt1=-2.3572041e-008 wkt1=-3.9150482e-007            pkt1=1.4774804e-014             kt2=0.060915125 wkt2=-1.0468272e-007            ute=-0.5                       ua1=-5.8438997e-009 lua1=1.3925378e-016             wua1=4.4893292e-015             pua1=-1.5789198e-022 ub1=5.7384557e-018             lub1=-8.939514e-026             wub1=-4.7846601e-024 pub1=1.663284e-031              uc1=-1.7193937e-010            luc1=4.114012e-018 wuc1=9.6606375e-017             puc1=-5.4369372e-025            at=-37221.966 lu0=2.0942689e-010             pu0=-1.860071e-016             lpdiblc2=5.0435e-010 wpdiblc2=4.80935e-009               ppdiblc2=-3.174171e-016             laigbinv=-2.5622263e-010 paigbinv=2.3213771e-016             lbigc=-1.2181825e-010            pbigc=8.1049877e-017 lbigsd=4.8353794e-011             pbigsd=-3.5229992e-017            lkt2=-3.2547331e-009 pkt2=3.5373637e-015             lat=0.0025491024               wat=0.042375329 pat=-1.5749003e-009            letab=1.5828692e-009             petab=4.1822708e-015 leta0=5.0876759e-009             weta0=-1.0362431e-008            peta0=3.154827e-016 lvsat=-0.00016492358             pvsat=7.6029096e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' voff_ff=-0.0184556                 voff_ss=0.0276833                  voff_mcl=-0.0256666 lvoff_ff=7.75133e-10                lvoff_ss=-1.1627e-09                lvoff_mcl=1.078e-09 wvoff_ff=1.00767e-08                wvoff_ss=-1.51151e-08               wvoff_mcl=3.3e-14 pvoff_ff=-4.23223e-16               pvoff_ss=6.34834e-16                pvoff_mcl=-2e-22 u0_ff=0.000461389                u0_ss=-0.000461389               wu0_ff=-2.51918e-10 wu0_ss=2.51918e-10                vsat_ff=3097.22                    vsat_ss=1516.67 vsat_sf=-886.113                   vsat_fs=10113.9                    wvsat_ff=-0.00114508 wvsat_ss=-0.0013741                 wvsat_sf=-0.00251918                wvsat_fs=-0.00251915 ua1_ff=2.78056e-10                ua1_sf=1.11222e-10                ua1_fs=-1.11222e-10 ua1_ss=-5.12945e-10               lua1_ff=-1.16783e-17               lua1_sf=-4.67133e-18 lua1_fs=4.67133e-18                lua1_ss=1.94297e-17                wua1_ff=-2.51918e-16 wua1_sf=-1.00767e-16               wua1_fs=1.00767e-16                wua1_ss=3.80167e-16 pua1_ff=1.05806e-23                pua1_sf=4.23223e-24                pua1_fs=-4.23223e-24 pua1_ss=-1.48128e-23               lu0_ff=-1.93783e-11               lu0_ss=1.93783e-11 pu0_ff=1.05806e-17                pu0_ss=-1.05806e-17               lvsat_ff=-0.000193783 lvsat_ss=3.3e-10                    lvsat_sf=3.7217e-05                 lvsat_fs=-0.000424783 pvsat_ff=1.05806e-10                pvsat_ss=4e-16                      pvsat_sf=1.05806e-10 pvsat_fs=1.05806e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.15 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.4854928 lvth0=2.3930385e-008             wvth0=-4.5172086e-010            pvth0=-1.9685274e-015 k2=-0.0029478821              lk2=9.2782448e-009             wk2=-2.9631107e-009 pk2=-7.6846549e-016            cit=0.0016721264               lcit=-4.1658957e-014 wcit=-2.424918e-010             pcit=1.1566619e-020             voff=-0.14565146 lvoff=-6.9056162e-012            wvoff=-6.9794208e-010            pvoff=2.4779257e-018 eta0=0.12436489                 etab=-0.20372022                wetab=1.7586781e-008 u0=0.010552524                wu0=-2.3670435e-010            ua=1.9187061e-010 lua=-2.5571457e-016            wua=-9.3130185e-017            pua=2.826312e-023 ub=1.0776882e-018             lub=3.5142448e-026             wub=-9.1201228e-027 pub=-7.3810323e-033            uc=-5.4008815e-010            luc=3.6067307e-016 wuc=5.5627289e-018             puc=-5.0047872e-023            vsat=95111.111 wvsat=-0.0027906667              a0=2.1500748                  la0=-2.7602892e-012 wa0=-1.8019343e-007            pa0=7.6183983e-019             ags=1.0489911 lags=6.229998e-007              wags=-1.5744241e-007            pags=-9.3774562e-014 keta=-0.25907647                lketa=2.8196155e-007             wketa=3.2399987e-008 pketa=-3.7351978e-014            pclm=0.17860212                 lpclm=6.9309452e-012 wpclm=-9.1141047e-009            ppclm=-1.9129409e-018            pdiblc2=0.0005 aigbacc=0.012678585                laigbacc=-7.2093943e-011            waigbacc=-2.5029869e-010 paigbacc=9.9039734e-018             aigbinv=0.010967067                waigbinv=-5.19064e-011 aigc=0.0062199203               laigc=1.9554155e-011             waigc=-8.487808e-011 paigc=-4.946626e-018             bigc=0.0017035178               wbigc=-1.0091051e-010 aigsd=0.0046761536               laigsd=5.2055128e-011             waigsd=1.4689984e-010 paigsd=-2.8421469e-017            bigsd=1.9872222e-005             wbigsd=7.8557267e-011 tvoff=0.00255474                 ltvoff=-8.33271e-010              wtvoff=-5.52911e-011 ptvoff=3.99935e-017               kt1=-0.2532411                 lkt1=-3.0548582e-009 wkt1=3.2327638e-008             pkt1=-8.8115006e-015            kt2=-0.088444444 wkt2=1.1162667e-008             ute=-1.4819409                 wute=1.4318352e-007 ua1=3.9676144e-009             lua1=-1.0223332e-017            wua1=-1.0746777e-015 pua1=5.5809272e-024             ub1=-6.2898419e-018            lub1=8.2659891e-030 wub1=1.8178204e-024             pub1=-2.3372356e-036            uc1=9.0666568e-010 luc1=-8.4155052e-016            wuc1=2.3950683e-016             puc1=-1.9544368e-022 at=100000                     lu0=0                          pu0=0 lat=0                          wat=0                          pat=0 leta0=0                          weta0=-2.3832293e-009            peta0=0 lvsat=0                          pvsat=0                          jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)' jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                ua1_ff=1.11833e-11 ua1_ss=-1.11833e-11               ua1_fs=-1.11833e-11               ua1_sf=1.11833e-11 lua1_ff=-1.00728e-16               lua1_ss=1.00728e-16                lua1_fs=1.00728e-16 lua1_sf=-1.00728e-16               wua1_ff=-3.08659e-18               wua1_ss=3.08659e-18 wua1_fs=3.08659e-18                wua1_sf=-3.08659e-18               pua1_ff=2.7801e-23 pua1_ss=-2.7801e-23                pua1_fs=-2.7801e-23                pua1_sf=2.7801e-23 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.16 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.4632581 lvth0=3.9858572e-009             wvth0=-3.0633178e-009            pvth0=3.740751e-016 k2=0.0094116987               lk2=-1.8082991e-009            wk2=-2.9100869e-009 pk2=-8.1602791e-016            cit=0.0016777626               lcit=-5.0972532e-012 wcit=-3.1599344e-010            pcit=6.5942538e-017             voff=-0.14148476 lvoff=-3.7444313e-009            wvoff=-1.7193674e-009            pvoff=9.1869639e-016 eta0=0.12436489                 etab=-0.20372022                wetab=1.7586781e-008 u0=0.010808022                wu0=-5.1396601e-010            ua=4.6137422e-010 lua=-4.974593e-016             wua=-1.6058779e-016            pua=8.8772591e-023 ub=9.4996548e-019             lub=1.4970977e-025             wub=1.4982734e-026 pub=-2.9001295e-032            uc=-1.551935e-010             luc=1.5422566e-017 wuc=-4.6267951e-017            puc=-3.5557519e-024            vsat=95111.111 wvsat=-0.0027906667              a0=3.1455925                  la0=-8.9298218e-007 wa0=-5.0943414e-007            pa0=2.9532968e-013             ags=2.6672978 lags=-8.2862132e-007            wags=-7.3018363e-007            pags=4.1997431e-013 keta=0.057335506                lketa=-1.8599944e-009            wketa=-6.5837147e-009 pketa=-2.3835971e-015            pclm=0.047936114                lpclm=1.1721434e-007 wpclm=-2.0783483e-009            ppclm=-6.3129864e-015            pdiblc2=0.0001016485 aigbacc=0.013610585                laigbacc=-9.080982e-010             waigbacc=-4.134762e-010 paigbacc=1.562742e-016              aigbinv=0.013776169                waigbinv=-1.0986371e-009 aigc=0.0071675701               laigc=-8.3048773e-010            waigc=-4.6196379e-010 paigc=3.3329925e-016             bigc=0.0028104002               wbigc=-5.3529266e-010 aigsd=0.0042826868               laigsd=4.0499482e-010             waigsd=2.6955759e-010 paigsd=-1.3844547e-016            bigsd=-0.00047508922             wbigsd=2.4779166e-010 tvoff=0.00203183                 ltvoff=-3.64217e-010              wtvoff=-1.52161e-010 ptvoff=1.26886e-016               kt1=-0.21790575                lkt1=-3.4750662e-008 wkt1=1.1952109e-008             pkt1=9.4653495e-015             kt2=-0.10558184 wkt2=1.4428379e-008             ute=-1.8140992                 wute=2.4915392e-007 ua1=3.03934e-009               lua1=8.224388e-016              wua1=-6.5501423e-016 pua1=-3.708572e-022             ub1=-6.0610111e-018            lub1=-2.0525296e-025 wub1=1.4990462e-024             pub1=2.8593814e-031             uc1=3.9039959e-010 luc1=-3.7845984e-016            wuc1=-1.4025915e-016            puc1=1.4520641e-022 at=42988.026                  lu0=-2.2918223e-010            pu0=2.4870371e-016 lpdiblc2=3.573213e-010              wpdiblc2=-4.7963607e-010            ppdiblc2=4.3023355e-016 laigbinv=-2.519765e-009             paigbinv=9.3891743e-016             lbigc=-9.9287349e-010 pbigc=3.8964079e-016             lbigsd=4.4398042e-010             pbigsd=-1.5180326e-016 lkt2=1.5372244e-008             pkt2=-2.9293438e-015            lute=2.97946e-007 pute=-9.5055444e-014            lat=0.051139741                wat=0.031128538 pat=-2.7922298e-008            leta0=0                          weta0=-2.3832293e-009 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' ua1_ff=-2.01548e-10               ua1_ss=2.01548e-10                ua1_fs=2.01548e-10 ua1_sf=-1.01111e-10               lua1_ff=9.0092e-17                 lua1_ss=-9.0092e-17 lua1_fs=-9.0092e-17                lua1_sf=-2.2e-23                   wua1_ff=5.56273e-17 wua1_ss=-5.56273e-17               wua1_fs=-5.56273e-17               wua1_sf=2.79067e-17 pua1_ff=-2.48654e-23               pua1_ss=2.48654e-23                pua1_fs=2.48654e-23 pua1_sf=-2e-30 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.17 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.46813694 lvth0=6.1666995e-009             wvth0=-3.1141364e-009            pvth0=3.9679095e-016 k2=0.013446521                lk2=-3.6118647e-009            wk2=-6.7878945e-009 pk2=9.1735211e-016             cit=0.00079652947              lcit=3.8881394e-010 wcit=-4.3613778e-011            pcit=-5.5811171e-017            voff=-0.14944454 lvoff=-1.8640863e-010            wvoff=1.1862035e-009             pvoff=-3.8009376e-016 eta0=0.12436489                 etab=-0.20372022                wetab=1.7586781e-008 u0=0.0098517737               wu0=2.5427267e-010             ua=-1.1156897e-010 lua=-2.413537e-016             wua=8.5777481e-017             pua=-2.1352684e-023 ub=1.3071612e-018             lub=-9.9567125e-027            wub=-1.2051794e-025 pub=3.1567506e-032             uc=-8.5314501e-011            luc=-1.5813344e-017 wuc=-9.3418282e-017            puc=1.7520446e-023             vsat=91355.23 wvsat=-0.00073995543             a0=1.2371592                  la0=-3.9912506e-008 wa0=3.2638722e-007             pa0=-7.828247e-014             ags=1.2527777 lags=-1.9633087e-007            wags=2.82106e-007               pags=-3.2519156e-014 keta=0.043417993                lketa=4.361134e-009              wketa=-5.918174e-009 pketa=-2.6810938e-015            pclm=0.054751769                lpclm=1.1416774e-007 wpclm=-8.1407044e-009            ppclm=-3.6031132e-015            pdiblc2=-0.00068074122 aigbacc=0.012491991                laigbacc=-4.0808644e-010            waigbacc=-5.2750221e-010 paigbacc=2.0724383e-016             aigbinv=0.009144457                waigbinv=8.494868e-010 aigc=0.004655152                laigc=2.9256317e-010             waigc=4.9054861e-010 paigc=-9.2473787e-017            bigc=-0.00011406599             wbigc=5.6310102e-010 aigsd=0.0054367358               laigsd=-1.1086508e-010            waigsd=-1.1029399e-010 paigsd=3.1348188e-017             bigsd=0.00081655945              wbigsd=-1.6254796e-010 tvoff=0.00198205                 ltvoff=-3.41966e-010              wtvoff=-7.0291e-011 ptvoff=9.02898e-017               kt1=-0.25947675                lkt1=-1.6168427e-008 wkt1=2.4724197e-008             pkt1=3.7562258e-015             kt2=-0.090754943 wkt2=1.2917428e-008             ute=-1.0732744                 wute=2.5020116e-008 ua1=6.4650426e-009             lua1=-7.0885028e-016            wua1=-1.8335479e-015 pua1=1.5594735e-022             ub1=-8.5321528e-018            lub1=8.9934739e-025 wub1=2.5689809e-024             pub1=-1.9232266e-031            uc1=-5.0880443e-010 luc1=2.3484362e-017             wuc1=1.8577371e-016             puc1=-5.3028293e-025 at=132064.89                  lu0=1.9826131e-010             pu0=-9.4698976e-017 lpdiblc2=7.070495e-010              wpdiblc2=7.9755053e-010             ppdiblc2=-1.4066886e-016 laigbinv=-4.4938959e-010            paigbinv=6.810605e-017              lbigc=3.1436288e-010 pbigc=-1.0134119e-016            lbigsd=-1.3338654e-010            pbigsd=3.1618558e-017 lkt2=8.7446208e-009             pkt2=-2.2539488e-015            lute=-3.3202689e-008 pute=5.1323666e-015             lat=0.011322381                wat=-0.017507432 pat=-6.1820201e-009            leta0=0                          weta0=-2.3832293e-009 peta0=0                          lvsat=0.001678879                pvsat=-9.1666792e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' ua1_sf=-1.93148e-10               lua1_sf=4.11406e-17                wua1_sf=5.33089e-17 pua1_sf=-1.13548e-23 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.18 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.44001431 lvth0=1.7657917e-010             wvth0=-3.9041527e-009            pvth0=5.6506445e-016 k2=-0.005331372               lk2=3.8782651e-010             wk2=-1.3688674e-009 pk2=-2.3690066e-016            cit=0.0021049197               lcit=1.1012683e-010 wcit=-3.8143955e-010            pcit=1.6145719e-017             voff=-0.13047127 lvoff=-4.2277159e-009            wvoff=-2.675748e-009             pvoff=4.425019e-016 eta0=0.12436489                 etab=-0.20372022                wetab=1.7586781e-008 u0=0.011197167                wu0=-2.6211935e-010            ua=-9.7537449e-010 lua=-5.7363118e-017            wua=-5.2824883e-017            pua=8.1696193e-024 ub=1.189132e-018              lub=1.5183517e-026             wub=1.0828298e-025 pub=-1.716709e-032             uc=-2.3584995e-010            luc=1.6250707e-017 wuc=-9.162556e-018             puc=-4.2602357e-025            vsat=102086.32 wvsat=-0.0065991304              a0=3.0167232                  la0=-4.1895963e-007 wa0=-9.2150303e-008            pa0=1.0866023e-014             ags=-0.13086674 lags=9.8385407e-008             wags=2.1880494e-007             pags=-1.9036029e-014 keta=0.18220481                 lketa=-2.5200457e-008            wketa=-5.5381883e-008 pketa=7.8546762e-015             pclm=0.76319086                 lpclm=-3.6729786e-008 wpclm=-5.241056e-008             ppclm=5.8263661e-015             pdiblc2=0.0023892986 aigbacc=0.011189679                laigbacc=-1.3069406e-010            waigbacc=4.4386521e-010 paigbacc=3.4256728e-019             aigbinv=0.0050050932               waigbinv=1.9765614e-009 aigc=0.0059460145               laigc=1.7609463e-011             waigc=1.0479788e-010 paigc=-1.0308882e-017            bigc=0.0012423054               wbigc=1.5070109e-010 aigsd=0.0047311831               laigsd=3.9417639e-011             waigsd=5.9045466e-011 paigsd=-4.7211161e-018            bigsd=7.4123185e-005             wbigsd=4.4827409e-012 tvoff=0.00044093                 ltvoff=-1.37079e-011              wtvoff=4.16223e-010 ptvoff=-1.33378e-017              kt1=-0.35946409                lkt1=5.1288764e-009 wkt1=6.0990103e-008             pkt1=-3.968412e-015             kt2=-0.06539894 wkt2=1.1337615e-008             ute=-1.3433833                 wute=8.26436e-008 ua1=4.6619799e-009             lua1=-3.2479793e-016            wua1=-1.7023572e-015 pua1=1.2800373e-022             ub1=-6.3750778e-018            lub1=4.398904e-025 wub1=2.5478159e-024             pub1=-1.8781451e-031            uc1=-5.7806703e-010 luc1=3.8237296e-017             wuc1=2.6154705e-016             puc1=-1.6670003e-023 at=245494.23                  lu0=-8.8307569e-011            pu0=1.5292522e-017 lpdiblc2=5.3131024e-011             wpdiblc2=2.3182068e-010             ppdiblc2=-2.0168399e-017 laigbinv=4.3229489e-010             paigbinv=-1.7196084e-016            lbigc=2.5455765e-011 pbigc=-1.3499999e-017            lbigsd=2.4752383e-011             pbigsd=-3.9589821e-018 lkt2=3.3437923e-009             pkt2=-1.9174487e-015            lute=2.4330517e-008 pute=-7.1414356e-015            lat=-0.012838068               wat=-0.067780436 pat=4.5261299e-009             leta0=0                          weta0=-2.3832293e-009 peta0=0                          lvsat=-0.00060684312             pvsat=3.3133634e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=690.48                     wvsat_ff=-2.2e-10                   ua1_fs=-6.98148e-11 lua1_fs=1.48706e-17                wua1_fs=1.92689e-17                pua1_fs=-4.10427e-24 lvsat_ff=-0.000147071               pvsat_ff=3.3e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.19 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.41905981 lvth0=-1.6464626e-009            wvth0=-2.809036e-009             pvth0=4.6978929e-016 k2=0.032398828                lk2=-2.8947008e-009            wk2=-7.1515777e-009 pk2=2.6619514e-016             cit=0.0027586957               lcit=5.3248311e-011 wcit=-3.0623613e-010            pcit=9.603021e-018              voff=-0.14725671 lvoff=-2.7673829e-009            wvoff=8.1195888e-011             pvoff=2.0264778e-016 eta0=0.12842694                 etab=-0.32263868                wetab=5.0408277e-008 u0=0.0095624228               wu0=5.0799468e-010             ua=-2.1130117e-009 lua=4.1611322e-017             wua=1.4905644e-016             pua=-9.3940558e-024 ub=2.0443023e-018             lub=-5.9216303e-026            wub=-1.8127472e-025 pub=8.0244299e-033             uc=9.8548518e-012             luc=-5.1256114e-018 wuc=-2.6409939e-017            puc=1.0744988e-024             vsat=121099.46 wvsat=-0.0093619501              a0=4.4878661                  la0=-5.4694906e-007 wa0=-2.4943386e-007            pa0=2.4549693e-014             ags=1 lags=0                          wags=0                          pags=0 keta=-0.13599368                lketa=2.482811e-009              wketa=2.1142556e-009 pketa=2.8525122e-015             pclm=0.35231171                 lpclm=-9.8330035e-010 wpclm=-1.6769129e-009            ppclm=1.4125388e-015             pdiblc2=0.000875 aigbacc=0.0098561041               laigbacc=-1.4673044e-011            waigbacc=2.1877609e-010 paigbacc=1.9925321e-017             aigbinv=0.009974                   aigc=0.0065602355 laigc=-3.5827769e-011            waigc=-3.8296283e-011            paigc=2.14031e-018 bigc=0.0019666808               wbigc=-5.7641912e-011            aigsd=0.0052802438 laigsd=-8.3506355e-012            waigsd=-9.8559359e-011            paigsd=8.9905038e-018 bigsd=0.00052392041              wbigsd=-1.4959303e-010            tvoff=-0.000745369 ltvoff=8.95001e-011               wtvoff=5.36763e-010               ptvoff=-2.38247e-017 kt1=-0.36651232                lkt1=5.7420729e-009             wkt1=3.9063499e-008 pkt1=-2.0607975e-015            kt2=-0.001874602               wkt2=-1.8200218e-008 ute=-1.3924519                 wute=1.5513781e-007             ua1=2.2725186e-009 lua1=-1.169148e-016             wua1=-4.5745487e-016            pua1=1.969723e-023 ub1=-3.2258547e-018            lub1=1.6590799e-025             wub1=7.8653963e-025 pub1=-3.4583475e-032            uc1=-5.1778895e-010            luc1=3.2993103e-017 wuc1=1.7897492e-016             puc1=-9.486228e-024             at=158876.52 lu0=5.3915194e-011             pu0=-5.1707398e-017            lpdiblc2=1.84875e-010 lbigc=-3.7564896e-011            pbigc=4.6258417e-018             lbigsd=-1.4379975e-011 pbigsd=9.4456102e-018             lkt2=-2.1828251e-009            pkt2=6.5234278e-016 lute=2.8599478e-008             pute=-1.3448432e-014            lat=-0.0053023271 wat=-0.034244573               pat=1.6085098e-009             letab=1.0345906e-008 petab=-2.8554701e-015            leta0=-3.5339872e-010            weta0=5.9167347e-009 peta0=-7.2209687e-016            lvsat=-0.0022609862              pvsat=5.7170166e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=-2416.67                   wvsat_ff=-2.2e-09                   ua1_ff=-7.24074e-11 ua1_ss=-7.08336e-11               ua1_fs=1.73518e-10                lua1_ff=6.29944e-18 lua1_ss=6.16246e-18                lua1_fs=-6.2994e-18                wua1_ff=3.95344e-17 wua1_ss=-4.4e-23                   wua1_fs=-6.74411e-17               pua1_ff=-3.4395e-24 pua1_ss=-3.3e-30                   pua1_fs=3.4395e-24                 lvsat_ff=0.00012325 pvsat_ff=3.3e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.20 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.46438086 lvth0=6.649108e-010              wvth0=1.9032835e-008             pvth0=-6.4414611e-016 k2=0.021266859                lk2=-2.3269704e-009            wk2=1.0819374e-009 pk2=-1.5371414e-016            cit=-0.0026708067              lcit=3.3015293e-010 wcit=1.2078267e-009             pcit=-6.7614184e-017            voff=-0.16818969 lvoff=-1.6998009e-009            wvoff=7.141305e-009              pvoff=-1.5741778e-016 eta0=0.21658369                 etab=-0.2666383                 wetab=-5.5683102e-009 u0=0.015225818                wu0=-1.0811614e-009            ua=-1.2835537e-009 lua=-6.9103929e-019            wua=-5.2199941e-017            pua=8.7001959e-025 ub=1.5068787e-018             lub=-3.1807697e-026            wub=-1.7143465e-025 pub=7.5225863e-033             uc=-1.8803859e-010            luc=4.9669542e-018 wuc=-4.2213484e-018            puc=-5.7119365e-026            vsat=150428.53 wvsat=-0.02868437                a0=25.703278                  la0=-1.6289351e-006 wa0=-6.2390144e-006            pa0=3.300183e-013              ags=1 lags=0                          wags=0                          pags=0 keta=0.46138518                 lketa=-2.7983511e-008            wketa=-9.6743111e-009 pketa=3.4537291e-015             pclm=-0.35972488                lpclm=3.5330566e-008 wpclm=2.5216601e-007             ppclm=-1.1533451e-014            pdiblc2=0.016374074 aigbacc=-0.0052920331              laigbacc=7.5788195e-010             waigbacc=5.9053183e-009 paigbacc=-2.7008833e-016            aigbinv=0.009974                   aigc=0.0073431551 laigc=-7.5756665e-011            waigc=-4.1352856e-010            paigc=2.1277156e-017 bigc=0.0026512431               wbigc=-4.331271e-010             aigsd=0.004277944 laigsd=4.2766653e-011             waigsd=2.3333284e-010             paigsd=-7.9359986e-018 bigsd=-1.8343271e-005            wbigsd=6.8658387e-011             tvoff=-0.00543839 ltvoff=3.28844e-010               wtvoff=1.86475e-009               ptvoff=-9.15522e-017 kt1=-0.7818271                 lkt1=2.6923127e-008             wkt1=1.2015157e-007 pkt1=-6.1962891e-015            kt2=-0.031643927               wkt2=-1.3878176e-008 ute=-3.3335815                 wute=-9.4231511e-008            ua1=8.9767274e-009 lua1=-4.5882944e-016            wua1=-2.3310708e-015            pua1=1.1525164e-022 ub1=-1.5560881e-17             lub1=7.9499434e-25              wub1=3.8441811e-24 pub1=-1.9052319e-31             uc1=-8.8954526e-011            luc1=1.1122547e-017 wuc1=2.0637641e-016             puc1=-1.0883704e-023            at=288583.52 lu0=-2.3491796e-010            pu0=2.9339561e-017             lpdiblc2=-6.0557778e-010 wpdiblc2=-5.2092444e-009            ppdiblc2=2.6567147e-016             lbigc=-7.2477569e-011 pbigc=2.3775587e-017             lbigsd=1.3275472e-011             pbigsd=-1.6852122e-018 lkt2=-6.6458958e-010            pkt2=4.3191863e-016             lute=1.2759709e-007 pute=-7.3059653e-016            lat=-0.011917384               wat=-0.085573018 pat=4.2262605e-009             letab=7.4898864e-009             petab=-6.6417867e-019 leta0=-4.849393e-009             weta0=-3.1216941e-008            peta0=1.1717206e-015 lvsat=-0.003756769               pvsat=1.5571451e-009 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=-14207.4                   vsat_ss=9437.04                    wvsat_ff=0.00520924 wvsat_ss=-0.00260462                ua1_fs=7.60371e-10                ua1_ss=8.55778e-10 ua1_ff=5.11115e-11                ua1_sf=-2.38519e-10               lua1_fs=-3.62288e-17 lua1_ss=-4.10946e-17               lua1_ff=4.4e-23                    lua1_sf=1.21644e-17 wua1_fs=-2.60462e-16               wua1_ss=-3.12555e-16               wua1_ff=-2.79069e-17 wua1_sf=1.30231e-16                pua1_fs=1.32836e-23                pua1_ss=1.59403e-23 pua1_ff=3.3e-30                    pua1_sf=-6.64179e-24               lvsat_ff=0.000724578 lvsat_ss=-0.000481289               pvsat_ff=-2.65672e-10               pvsat_ss=1.32836e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.21 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.46152009 lvth0=5.4475855e-010             wvth0=2.0164515e-008             pvth0=-6.9167671e-016 k2=0.046649434                lk2=-3.3930386e-009            wk2=-1.5658446e-008 pk2=5.4938197e-016             cit=0.00073090416              lcit=1.8728108e-010 wcit=-9.5578763e-010            pcit=2.3257618e-017             voff=-0.18034276 lvoff=-1.1893719e-009            wvoff=1.4951691e-008             pvoff=-4.8545398e-016 eta0=-0.065349101               etab=-0.25768802                wetab=-3.3257627e-008 u0=0.01457247                 wu0=-1.3736151e-009            ua=-1.4721923e-009 lua=7.2317808e-018             wua=-1.6735963e-018            pua=-1.2520869e-024 ub=1.1232419e-018             lub=-1.5694953e-026            wub=-9.429637e-026 pub=4.2827786e-033             uc=-2.1009419e-010            luc=5.8932891e-018 wuc=2.0951395e-017             puc=-1.1143746e-024            vsat=-9932.0313 wvsat=0.031151225                a0=-20.487361                 la0=3.1107178e-007 wa0=9.4332902e-006             pa0=-3.2821849e-013            ags=1 lags=0                          wags=0                          pags=0 keta=0.1594963                  lketa=-1.5304178e-008            wketa=4.9822702e-007 pketa=-1.7878127e-014            pclm=0.3246368                  lpclm=6.5873748e-009 wpclm=4.3937181e-008             ppclm=-2.7878396e-015            pdiblc2=0.0019148148 aigbacc=0.019295043                laigbacc=-2.7477526e-010            waigbacc=-1.8037959e-009 paigbacc=5.3694462e-017             aigbinv=0.0018399482               waigbinv=2.2449983e-009 aigc=0.0042850179               laigc=5.2685095e-011             waigc=4.3971801e-010 paigc=-1.45592e-017              bigc=-0.00022915406             wbigc=4.1732494e-010 aigsd=0.0061886225               laigsd=-3.7481844e-011            waigsd=-7.4660324e-011 paigsd=4.9997145e-018             bigsd=0.00088467276              wbigsd=-8.1721325e-011 tvoff=0.00339842                 ltvoff=-4.23019e-011              wtvoff=-1.19983e-009 ptvoff=3.71605e-017               kt1=-0.06051573                lkt1=-3.3719511e-009 wkt1=-1.1655901e-007            pkt1=3.7455553e-015             kt2=-0.10542424 wkt2=-1.3861429e-008            ute=0.45407407                 wute=-5.2092444e-007 ua1=-1.7853607e-010            lua1=-7.4308378e-017            wua1=1.3960407e-015 pua1=-4.1287039e-023            ub1=1.5137215e-18              lub1=7.786103e-26 wub1=-2.4779553e-24             pub1=7.5006535e-32              uc1=4.4425461e-010 luc1=-1.1272236e-017            wuc1=-2.3983554e-016            puc1=7.8571979e-024 at=-71628.29                  lu0=-2.0747735e-010            pu0=4.1622618e-017 lpdiblc2=1.7111111e-012             wpdiblc2=2.1395111e-009             ppdiblc2=-4.2976267e-017 laigbinv=3.4163018e-010             paigbinv=-9.4289929e-017            lbigc=4.849911e-011 pbigc=-1.1943399e-017            lbigsd=-2.4651201e-011            pbigsd=4.6307357e-018 lkt2=2.4341836e-009             pkt2=4.3121526e-016             lute=-3.1484444e-008 pute=1.7190507e-014             lat=0.0032115119               wat=0.061161182 pat=-1.9365759e-009            letab=7.1139748e-009             petab=1.1622871e-015 leta0=6.9917844e-009             weta0=1.3923086e-008             peta0=-7.2416054e-016 lvsat=0.0029783747               pvsat=-9.559499e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vth0_ff=0.0074963                  lvth0_ff=-3.14844e-10               wvth0_ff=-4.09298e-09 pvth0_ff=1.71905e-16                voff_ss=-0.0074963                 voff_ff=0.0112444 voff_mcl=-0.033163                  lvoff_ss=3.14844e-10                lvoff_ff=-4.72267e-10 lvoff_mcl=1.39285e-09                wvoff_ss=4.09298e-09                wvoff_ff=-6.13947e-09 wvoff_mcl=4.09296e-09                pvoff_ss=-1.71905e-16               pvoff_ff=2.57858e-16 pvoff_mcl=-1.71905e-16               u0_ff=-0.000374815               u0_mc=0.00187407 wu0_ff=2.04649e-10                wu0_mc=-1.02324e-09               vsat_ff=4918.53 vsat_ss=-2022.23                   vsat_sf=-11122.2                   vsat_fs=11122.2 vsat_mc=-5622.22                   wvsat_ff=-0.00213951                wvsat_ss=0.000558132 wvsat_sf=0.00306973                 wvsat_fs=-0.00306973                wvsat_mc=0.00306973 a0_sf=1.49926                    la0_sf=-6.29689e-08               wa0_sf=-8.18596e-07 pa0_sf=3.4381e-14                 ua1_ff=-1.32222e-10               ua1_sf=9.02225e-11 ua1_fs=-3.28741e-10               ua1_ss=-2.01704e-10               lua1_ff=7.69999e-18 lua1_sf=-1.64267e-18               lua1_fs=9.51378e-18                lua1_ss=3.3196e-18 wua1_ff=-2.79071e-17               wua1_sf=-8.93013e-17               wua1_fs=2.19532e-16 wua1_ss=2.10231e-16                pua1_ff=-3.3e-30                   pua1_sf=2.57858e-24 pua1_fs=-6.87621e-24               pua1_ss=-6.01668e-24               lu0_ff=1.57422e-11 lu0_mc=-7.87111e-11               pu0_ff=-8.59525e-18               pu0_mc=4.29763e-17 lvsat_ff=-7.87114e-05               lvsat_ss=2.2e-10                    lvsat_sf=0.000467133 lvsat_fs=-0.000467133               lvsat_mc=0.000236133                pvsat_ff=4.2976e-11 pvsat_ss=-3.3e-17                   pvsat_sf=-1.28929e-10               pvsat_fs=1.28929e-10 pvsat_mc=-1.28929e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.22 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.48066923 lvth0=1.9086375e-008             wvth0=-1.7830273e-009            pvth0=-6.3158063e-016 k2=-0.021256562               lk2=6.6586024e-009             wk2=2.0900849e-009 pk2=-4.5444191e-017            cit=0.00094774753              lcit=1.9439592e-016 wcit=-4.2563219e-011            pcit=1.5093803e-023             voff=-0.15276127 lvoff=1.4673054e-012             wvoff=1.2643681e-009             pvoff=1.6699938e-019 eta0=0.1338363                  etab=-0.14703704                wetab=1.9422222e-009 u0=0.0090200051               wu0=1.8627101e-010             ua=-2.036705e-011 lua=-2.7443837e-016            wua=-3.4552589e-017            pua=3.3430889e-023 ub=9.29467e-019               lub=1.0905459e-026             wub=3.1788941e-026 pub=-6.9162319e-034            uc=-5.043476e-010             luc=3.9115352e-017 wuc=-4.3016626e-018            puc=3.8702058e-023             vsat=85000 wvsat=0                          a0=1.5197322                  la0=3.2462052e-012 wa0=-6.218896e-009             pa0=-8.9595264e-019            ags=0.5139946 lags=2.902659e-007              wags=-9.7833939e-009            pags=-1.9400061e-015 keta=-0.10299159                lketa=1.1893918e-007             wketa=-1.067944e-008 pketa=7.6421974e-015             pclm=0.10728444                 lpclm=0 wpclm=1.0569573e-008             ppclm=0                          pdiblc2=0.0005 aigbacc=0.011954137                laigbacc=-7.0212404e-011            waigbacc=-5.0351139e-011 paigbacc=9.3846685e-018             aigbinv=0.010994333                waigbinv=-5.9432e-011 aigc=0.0059359726               laigc=2.9639732e-013             waigc=-6.5085171e-012 paigc=3.6851519e-019             bigc=0.0013633741               wbigc=-7.0308444e-012 aigsd=0.0051996867               laigsd=-1.0777101e-010            waigsd=2.4047106e-012 paigsd=1.5690544e-017             bigsd=0.00032912963              wbigsd=-6.7977778e-012 tvoff=0.00186502                 ltvoff=-7.01969e-010              wtvoff=1.35072e-010 ptvoff=3.7541e-018                kt1=-0.16416341                lkt1=-4.9389312e-008 wkt1=7.7421968e-009             pkt1=3.9768087e-015             kt2=-0.048 ute=-1.0236504                 wute=1.6695342e-008             ua1=1.4104837e-009 lua1=3.1629191e-017             wua1=-3.6890964e-016            pua1=-5.9703691e-024 ub1=-1.6845572e-018            lub1=-3.7099805e-030            wub1=5.4676186e-025 pub1=9.6813198e-037             uc1=2.4064287e-009             luc1=-2.1840266e-015 wuc1=-1.7442776e-016            puc1=1.7507973e-022             at=156296.3 lu0=-2.4539348e-013            pu0=6.7728601e-020             lat=0 wat=-0.015537778               pat=0                          leta0=0 weta0=-4.9973378e-009            peta0=0                          lvsat=0 pvsat=0                          jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)' jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                ags_ff=-0.00778326 lags_ff=7.01038e-08                wags_ff=2.14818e-09                pags_ff=-1.93487e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.23 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.46741061 lvth0=7.1933946e-009             wvth0=-1.9172249e-009            pvth0=-5.1120538e-016 k2=-0.0066387629              lk2=-6.4535632e-009            wk2=1.5198405e-009 pk2=4.6606497e-016             cit=0.00040969801              lcit=4.8263062e-010 wcit=3.3992376e-011             pcit=-6.8670354e-017            voff=-0.15590069 lvoff=2.8175242e-009             wvoff=2.2594298e-009             pvoff=-8.9240334e-016 eta0=0.1338363                  etab=-0.14703704                wetab=1.9422222e-009 u0=0.0082934117               wu0=1.8006672e-010             ua=-2.0767576e-010 lua=-1.0642246e-016            wua=2.4070003e-017             pua=-1.9153576e-023 ub=1.1720603e-018             lub=-2.0670074e-025            wub=-4.631544e-026 pub=6.9368006e-032             uc=-3.7753807e-010            luc=-7.4632796e-017 wuc=1.5099151e-017             puc=2.1299528e-023             vsat=85000 wvsat=0                          a0=1.0799179                  la0=3.9451667e-007 wa0=6.0692037e-008             pa0=-6.0020003e-014            ags=-0.31928159 lags=1.0377146e-006             wags=9.4112273e-008             pags=-9.5134419e-014 keta=0.073544807                lketa=-3.9413973e-008            wketa=-1.1057482e-008 pketa=7.981301e-015              pclm=0.004990242                lpclm=9.17579e-008 wpclm=9.7747124e-009             ppclm=7.1299024e-016             pdiblc2=-0.0020908709 aigbacc=0.012490334                laigbacc=-5.5118054e-010            waigbacc=-1.0428677e-010 paigbacc=5.7764929e-017             aigbinv=0.0095279158               waigbinv=7.3880839e-011 aigc=0.0053767621               laigc=5.0190821e-010             waigc=3.2299222e-011 paigc=-3.4442027e-017            bigc=0.00075318044              wbigc=3.2499981e-011 aigsd=0.005184112                laigsd=-9.3800524e-011            waigsd=2.076424e-011 paigsd=-7.7795369e-019            bigsd=0.00043021049              wbigsd=-2.0710563e-012 tvoff=0.000828334                ltvoff=2.27937e-010               wtvoff=1.80003e-010 ptvoff=-3.65487e-017              kt1=-0.22585842                lkt1=5.9511133e-009 wkt1=1.4147045e-008             pkt1=-1.7683404e-015            kt2=-0.057038328 wkt2=1.0303693e-009             ute=-0.90319399                wute=-2.255917e-009 ua1=2.5746538e-009             lua1=-1.0126314e-015            wua1=-5.2676085e-016 pua1=1.3562217e-022             ub1=-3.4423858e-018            lub1=1.5767685e-024 wub1=7.7630562e-025             pub1=-2.0589978e-031            uc1=-2.9711726e-010 luc1=2.410541e-016              wuc1=4.9495505e-017             puc1=-2.577944e-023 at=251316.25                  lu0=6.5150887e-010             pu0=5.632969e-018 lpdiblc2=2.3240112e-009             wpdiblc2=1.2549928e-010             ppdiblc2=-1.1257285e-016 laigbinv=1.3153765e-009             paigbinv=-1.1958162e-016            lbigc=5.4734369e-010 pbigc=-3.5459151e-017            lbigsd=-9.0669535e-011            pbigsd=-4.2398692e-018 lkt2=8.1073798e-009             pkt2=-9.2424129e-016            lute=-1.0804938e-007 pute=1.6999279e-014             lat=-0.085232901               wat=-0.026370053 pat=9.7165507e-009             leta0=0                          weta0=-4.9973378e-009 peta0=0                          lvsat=0                          pvsat=0 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' u0_ff=-0.000174753               u0_sf=-0.000174753               wu0_ff=4.82319e-11 wu0_sf=4.82319e-11                ags_ff=0.140272                   lags_ff=-6.27014e-08 wags_ff=-3.8715e-08                pags_ff=1.73056e-14                lu0_ff=1.56754e-10 lu0_sf=1.56754e-10                pu0_ff=-4.3264e-17                pu0_sf=-4.3264e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.24 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.4712115 lvth0=8.8923858e-009             wvth0=-2.2655625e-009            pvth0=-3.5549845e-016 k2=-0.02485978                lk2=1.6912317e-009             wk2=3.7846447e-009 pk2=-5.4630249e-016            cit=0.00085443032              lcit=2.8383527e-010 wcit=-5.9594414e-011            pcit=-2.6837058e-017            voff=-0.14266936 lvoff=-3.0968812e-009            wvoff=-6.8374693e-010            pvoff=4.2319666e-016 eta0=0.1338363                  etab=-0.14703704                wetab=1.9422222e-009 u0=0.010336962                wu0=1.203605e-010              ua=3.8254643e-010 lua=-3.7025178e-016            wua=-5.0598369e-017            pua=1.4223186e-023 ub=2.5638787e-019             lub=2.0260484e-025             wub=1.694955e-025 pub=-2.7099482e-032            uc=-7.8528949e-010            luc=1.0763209e-016 wuc=9.9774814e-017             puc=-1.6550494e-023            vsat=90388.653 wvsat=-0.00047318031             a0=2.8971796                  la0=-4.177993e-007 wa0=-1.3177841e-007            pa0=2.6014285e-014             ags=3.0883641 lags=-4.8550297e-007            wags=-2.2451584e-007            pags=4.7292346e-014 keta=0.0057727901               lketa=-9.1198816e-009            wketa=4.4719019e-009 pketa=1.0396665e-015             pclm=-0.16052687                lpclm=1.6574405e-007 wpclm=5.12762e-008               ppclm=-1.7838175e-014            pdiblc2=0.0032602411 aigbacc=0.0096835307               laigbacc=7.0346036e-010             waigbacc=2.4763274e-010 paigbacc=-9.9543089e-017            aigbinv=0.013456071                waigbinv=-3.4051876e-010 aigc=0.0064919643               laigc=3.4128401e-012             waigc=-1.6411589e-011 paigc=-1.2668294e-017            bigc=0.0019859663               wbigc=-1.6507888e-011 aigsd=0.0051039234               laigsd=-5.79562e-011              waigsd=-1.8437751e-011 paigsd=1.6745336e-017             bigsd=0.0004426096               wbigsd=-5.9337802e-011 tvoff=0.00126667                 ltvoff=3.20002e-011               wtvoff=1.27153e-010 ptvoff=-1.2925e-017               kt1=-0.22271942                lkt1=4.5479778e-009 wkt1=1.4579174e-008             pkt1=-1.961502e-015             kt2=-0.041104544 wkt2=-7.8608202e-010            ute=-1.1464232                 wute=4.5209181e-008 ua1=1.2663249e-009             lua1=-4.2780836e-016            wua1=-3.9870182e-016 pua1=7.8379781e-023             ub1=-1.1528971e-018            lub1=5.5336707e-025 wub1=5.3230631e-025             pub1=-9.6832091e-032            uc1=1.1976644e-010 luc1=5.4707083e-017             wuc1=1.2288155e-017             puc1=-9.147754e-024 at=102854.81                  lu0=-2.6195835e-010            pu0=3.2321648e-017 lpdiblc2=-6.7935867e-011            wpdiblc2=-2.9016058e-010            ppdiblc2=7.3227104e-017 laigbinv=-4.4050898e-010            paigbinv=6.5655003e-017             lbigc=-3.7115894e-012 pbigc=-1.3552633e-017            lbigsd=-9.6211936e-011            pbigsd=2.1358366e-017 lkt2=9.8497841e-010             pkt2=-1.1228754e-016            lute=6.7407218e-010 pute=-4.2176194e-015            lat=-0.018870635               wat=-0.0094454481 pat=2.1512524e-009             leta0=0                          weta0=-4.9973378e-009 peta0=0                          lvsat=-0.002408728               pvsat=2.115116e-010 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' u0_ff=0.000143899                u0_sf=0.000143899                wu0_ff=-3.9716e-11 wu0_sf=-3.9716e-11                vsat_ff=-1281.1                    wvsat_ff=0.000353584 lu0_ff=1.43163e-11                lu0_sf=1.43163e-11                pu0_ff=-3.95131e-18 pu0_sf=-3.95131e-18               lvsat_ff=0.000572652                pvsat_ff=-1.58052e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.25 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.43371066 lvth0=9.0470953e-010             wvth0=-5.6439612e-009            pvth0=3.6410048e-016 k2=-0.016968441               lk2=1.037628e-011              wk2=1.8429635e-009 pk2=-1.327244e-016             cit=0.0016003348               lcit=1.2495761e-010 wcit=-2.4217413e-010            pcit=1.2052422e-017             voff=-0.14127037 lvoff=-3.3948666e-009            wvoff=3.0480317e-010             pvoff=2.1263549e-016 eta0=0.1338363                  etab=-0.14703704                wetab=1.9422222e-009 u0=0.0087399593               wu0=4.1607007e-010             ua=-1.3325399e-009 lua=-4.9383907e-018            wua=4.5752765e-017             pua=-6.2996056e-024 ub=1.4467454e-018             lub=-5.0941308e-026            wub=3.7181678e-026 pub=1.0833613e-033             uc=-4.1376124e-010            luc=2.8496571e-017 wuc=3.9940958e-017             puc=-3.8058821e-024            vsat=74992.501 wvsat=0.00087876344              a0=2.8532872                  la0=-4.0845022e-007 wa0=-4.704197e-008             pa0=7.9654242e-015             ags=0.67713157 lags=2.8089553e-008             wags=-4.2025989e-009            pags=3.6562611e-016 keta=-0.088373453               lketa=1.0933268e-008             wketa=1.9297716e-008 pketa=-2.118232e-015             pclm=0.81441966                 lpclm=-4.1919562e-008 wpclm=-6.6549711e-008            ppclm=7.2587442e-015             pdiblc2=0.0029007578 aigbacc=0.014326526                laigbacc=-2.8549759e-010            waigbacc=-4.219045e-010 paigbacc=4.3068342e-017             aigbinv=0.012509537                waigbinv=-9.4665038e-011 aigc=0.0066441398               laigc=-2.9000535e-011            waigc=-8.7884695e-011 paigc=2.5554771e-018             bigc=0.0021268674               wbigc=-9.3438007e-011 aigsd=0.0046767238               laigsd=3.3037308e-011             waigsd=7.4076243e-011 paigsd=-2.9601447e-018            bigsd=-7.5877435e-005            wbigsd=4.5882912e-011 tvoff=0.00159109                 ltvoff=-3.71002e-011              wtvoff=9.87801e-011 ptvoff=-6.88149e-018              kt1=-0.14772987                lkt1=-1.1424796e-008 wkt1=2.5514581e-009             pkt1=6.0040149e-016             kt2=-0.0096009212 wkt2=-4.0626378e-009            ute=-1.2589                    wute=5.9326195e-008 ua1=-2.1454089e-009            lua1=2.9889095e-016             wua1=1.7648212e-016 pua1=-4.4134398e-023            ub1=3.7072974e-018             lub1=-4.8185436e-025 wub1=-2.3491968e-025            pub1=6.6587046e-032             uc1=5.9015371e-010 luc1=-4.5485405e-017            wuc1=-6.0881873e-017            puc1=6.4374619e-024 at=-23446.848                 lu0=7.8203347e-011             pu0=-3.0664491e-017 lpdiblc2=8.6340733e-012             wpdiblc2=9.0657939e-011             ppdiblc2=-7.8872407e-018 laigbinv=-2.3889715e-010            paigbinv=1.3288161e-017             lbigc=-3.3723516e-011 pbigc=2.8334824e-018             lbigsd=1.4225803e-011             pbigsd=-1.0536459e-018 lkt2=-5.7252932e-009            pkt2=5.8561885e-016             lute=2.4631632e-008 pute=-7.2245434e-015            lat=0.0080316176               wat=0.0064473017 pat=-1.2339033e-009            leta0=0                          weta0=-4.9973378e-009 peta0=0                          lvsat=0.0008706524               pvsat=-7.6452419e-011 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' u0_ff=0.000211111                u0_sf=0.000211111                wu0_ff=-5.82667e-11 wu0_sf=-5.82667e-11               vsat_ff=3555.56                    wvsat_ff=-0.000790762 lu0_ff=1.3e-17                    lu0_sf=1.3e-17                    pu0_ff=-1.9e-24 pu0_sf=-1.9e-24                   lvsat_ff=-0.000457555               pvsat_ff=8.56936e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.26 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.41727114 lvth0=-5.2552815e-010            wvth0=-3.3027073e-009            pvth0=1.6041138e-016 k2=0.0090013032               lk2=-2.2489914e-009            wk2=-6.9386103e-010 pk2=8.7979337e-017             cit=0.002022501                lcit=8.8229159e-011 wcit=-1.0304638e-010            pcit=-5.1693153e-020            voff=-0.15390815 lvoff=-2.2953791e-009            wvoff=1.9169959e-009             pvoff=7.2374723e-017 eta0=0.18474717                 etab=-0.15261975                wetab=3.4830518e-009 u0=0.011384591                wu0=5.076257e-012              ua=-1.2715144e-009 lua=-1.0247612e-017            wua=-8.3196839e-017            pua=4.9190099e-024 ub=8.7371249e-019             lub=-1.0874466e-027            wub=1.4180807e-025 pub=-8.0191344e-033            uc=-7.7122068e-011            luc=-7.9103676e-019 wuc=-2.4043093e-018            puc=-1.2184385e-025            vsat=87530.705 wvsat=-9.6974259e-005            a0=2.0887495                  la0=-3.4193543e-007 wa0=4.1272231e-007             pa0=-3.2034068e-014            ags=1 lags=0                          wags=0                          pags=0 keta=-0.023554784               lketa=5.294044e-009              wketa=-2.891888e-008 pketa=2.0766119e-015             pclm=0.19986728                 lpclm=1.1546495e-008 wpclm=4.0397748e-008             ppclm=-2.0456847e-015            pdiblc2=0.00037654321 aigbacc=0.009445871                laigbacc=1.3911937e-010             waigbacc=3.3200042e-010 paigbacc=-2.2521386e-017            aigbinv=0.0097635926               waigbinv=5.8072444e-011 aigc=0.0067525485               laigc=-3.8432098e-011            waigc=-9.1374668e-011 paigc=2.8591048e-018             bigc=0.0020993548               wbigc=-9.4259917e-011 aigsd=0.0044845362               laigsd=4.9757626e-011             waigsd=1.2105592e-010 paigsd=-7.0473762e-018            bigsd=-0.00046382811             wbigsd=1.2302556e-010 tvoff=0.00161                    ltvoff=-3.8746e-011               wtvoff=-1.1332e-010 ptvoff=1.15712e-017               kt1=-0.22539245                lkt1=-4.6681509e-009 wkt1=1.1441429e-010             pkt1=8.124243e-016              kt2=-0.074960545 wkt2=1.9715021e-009             ute=-0.34121447                wute=-1.3500371e-007 ua1=1.7728488e-009             lua1=-4.1997467e-017            wua1=-3.19546e-016 pua1=-9.7995223e-025            ub1=-2.0298119e-018            lub1=1.7274148e-026 wub1=4.5643182e-025             pub1=6.4394656e-033             uc1=1.4481236e-010 luc1=-6.7407072e-018            wuc1=-3.9030415e-018            puc1=1.4803036e-024 at=83651.278                  lu0=-1.5187962e-010            pu0=5.091972e-018 lpdiblc2=2.2824074e-010             wpdiblc2=1.3757407e-010             ppdiblc2=-1.1968944e-017 lbigc=-3.1329921e-011            pbigc=2.9049885e-018             lbigsd=4.7977512e-011 pbigsd=-7.7650562e-018            lkt2=-3.9005911e-011            pkt2=6.0648674e-017 lute=-5.5207007e-008            pute=9.6821579e-015             lat=-0.0012859194 wat=-0.013482406               pat=4.9998126e-010             letab=4.856963e-010 petab=-1.3405218e-016            leta0=-4.4292457e-009            weta0=-9.6276469e-009 peta0=4.028369e-016              lvsat=-0.00022017131             pvsat=8.4367605e-012 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' u0_ff=0.000510185                u0_sf=0.000510185                wu0_ff=-1.40811e-10 wu0_sf=-1.40811e-10               vsat_ff=-4117.28                   wvsat_ff=0.00046937 ua1_ff=1.70525e-10                ua1_sf=4.98457e-11                ua1_fs=-1.40617e-10 ua1_ss=-1.20679e-10               lua1_ff=-1.48356e-17               lua1_sf=-4.33657e-18 lua1_fs=1.22337e-17                lua1_ss=1.04991e-17                wua1_ff=-2.75148e-17 wua1_sf=-1.37574e-17               wua1_fs=1.92604e-17                wua1_ss=1.37574e-17 pua1_ff=2.39378e-24                pua1_sf=1.19689e-24                pua1_fs=-1.67565e-24 pua1_ss=-1.19689e-24               lu0_ff=-2.60194e-11               lu0_sf=-2.60194e-11 pu0_ff=7.18137e-18                pu0_sf=7.18137e-18                lvsat_ff=0.000209981 pvsat_ff=-2.39379e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.27 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.40138259 lvth0=-1.3358445e-009            wvth0=1.645313e-009              pvth0=-9.1937652e-017 k2=0.025762322                lk2=-3.1038034e-009            wk2=-1.5881055e-010 pk2=6.0691763e-017             cit=0.00091814779              lcit=1.4455117e-010 wcit=2.1727527e-010             pcit=-1.6388097e-017            voff=-0.17781273 lvoff=-1.076246e-009             wvoff=9.7972636e-009             pvoff=-3.2951893e-016 eta0=0.044765924                etab=-0.27631407                wetab=-2.8977956e-009 u0=0.012075269                wu0=-2.1160971e-010            ua=-1.3991627e-009 lua=-3.7375486e-018            wua=-2.0291863e-017            pua=1.7108562e-024 ub=8.7457094e-019             lub=-1.1312277e-027            wub=3.0822795e-027 pub=-9.4411932e-034            uc=-2.3627605e-010            luc=7.3258163e-018 wuc=9.0921896e-018             puc=-7.081653e-025             vsat=43738.156 wvsat=0.00076217407              a0=4.9476634                  la0=-4.8774005e-007 wa0=-5.1046478e-007            pa0=1.5048473e-014             ags=1 lags=0                          wags=0                          pags=0 keta=0.18408333                 lketa=-5.2955e-009               wketa=6.6861e-008 pketa=-2.808162e-015             pclm=0.90049265                 lpclm=-2.4185399e-008 wpclm=-9.5654024e-008            ppclm=4.8929557e-015             pdiblc2=-0.0070740741 aigbacc=0.018012956                laigbacc=-2.9780195e-010            waigbacc=-5.2685858e-010 paigbacc=2.1280423e-017             aigbinv=0.0087816914               waigbinv=3.2907718e-010 aigc=0.0059336077               laigc=3.3338826e-012             waigc=-2.4493495e-011 paigc=-5.5183503e-019            bigc=0.0011843277               wbigc=-2.8258468e-011 aigsd=0.0055288739               laigsd=-3.5035948e-012            waigsd=-1.1192381e-010 paigsd=4.8345899e-018             bigsd=0.00083507805              wbigsd=-1.668859e-010 tvoff=0.000682977                ltvoff=8.53231e-012               wtvoff=1.75255e-010 ptvoff=-3.1461e-018               kt1=-0.40525461                lkt1=4.5048193e-009 wkt1=1.6217563e-008             pkt1=-8.8363035e-018            kt2=-0.11893765 wkt2=1.0214892e-008             ute=-4.1442038                 wute=1.2950026e-007 ua1=8.3215503e-010             lua1=5.9779149e-018             wua1=-8.3168827e-017 pua1=-1.3035188e-023            ub1=-2.445104e-18              lub1=3.8454043e-26 wub1=2.2422659e-25              pub1=1.8281932e-32              uc1=1.0281294e-009 luc1=-5.1789875e-017            wuc1=-1.0193875e-016            puc1=6.4801246e-024 at=-43065.428                 lu0=-1.8710417e-010            pu0=1.6142956e-017 lpdiblc2=6.0822222e-010             wpdiblc2=1.2624444e-009             ppdiblc2=-6.9337333e-017 laigbinv=5.0076963e-011             paigbinv=-1.3821242e-017            lbigc=1.5336459e-011 pbigc=-4.6108541e-019            lbigsd=-1.8266703e-011            pbigsd=7.0204281e-018 lkt2=2.2038266e-009             pkt2=-3.5976423e-016            lute=1.3874545e-007 pute=-3.8075441e-015            lat=0.0051766327               wat=0.0059620929 pat=-4.9168818e-010            letab=6.7941067e-009             petab=1.9137104e-016 leta0=2.7097977e-009             weta0=1.6204764e-008             peta0=-9.1461604e-016 lvsat=0.0020132487               pvsat=-3.5379804e-011 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vsat_ff=7950.62                    wvsat_ff=-0.00090637                a0_fs=-0.65679 la0_fs=3.34963e-08                wa0_fs=1.81274e-07                pa0_fs=-9.24498e-15 ua1_ff=-2.84568e-10               ua1_sf=3.62345e-10                ua1_fs=-2.32593e-10 ua1_ss=-4.71358e-10               lua1_ff=8.37403e-18                lua1_sf=-2.02741e-17 lua1_fs=1.69244e-17                lua1_ss=2.83837e-17                wua1_ff=6.47405e-17 wua1_sf=-3.56074e-17               wua1_fs=1.35955e-17                wua1_ss=5.37348e-17 pua1_ff=-2.31124e-24               pua1_sf=2.31125e-24                pua1_fs=-1.38675e-24 pua1_ss=-3.23574e-24               lvsat_ff=-0.000405481               pvsat_ff=4.62249e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_hvt_mac.28 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.39192487 lvth0=-1.733069e-009             wvth0=9.5623275e-010             pvth0=-6.2996284e-017 k2=0.0033115825               lk2=-2.1608723e-009            wk2=-3.6971989e-009 pk2=2.0930407e-016             cit=-0.0027530469              lcit=2.9874135e-010 wcit=5.7828683e-012             pcit=-7.5054163e-018            voff=-0.13361255 lvoff=-2.9326533e-009            wvoff=2.054154e-009              pvoff=-4.3083282e-018 eta0=-0.025716749               etab=-0.4264659                 wetab=1.3325069e-008 u0=0.0092098433               wu0=1.0646996e-010             ua=-1.5147892e-009 lua=1.1187681e-018             wua=1.0083174e-017             pua=4.351046e-025 ub=7.5140066e-019             lub=4.0419239e-027             wub=8.3318044e-027 pub=-1.1645994e-033            uc=-4.2728272e-012            luc=-2.418319e-018 wuc=-3.58553e-017              puc=1.1796293e-024             vsat=99350.413 wvsat=0.00098926883              a0=19.381355                  la0=-1.0939551e-006 wa0=-1.5704754e-006            pa0=5.9568921e-014             ags=1 lags=0                          wags=0                          pags=0 keta=2.333642                   lketa=-9.5576963e-008            wketa=-1.0183718e-007 pketa=4.2771618e-015             pclm=0.67912943                 lpclm=-1.4888144e-008 wpclm=-5.3902783e-008            ppclm=3.1394036e-015             pdiblc2=0.013654321 aigbacc=0.015424294                laigbacc=-1.8907814e-010            waigbacc=-7.3546893e-010 paigbacc=3.0042058e-017             aigbinv=0.009974                   aigc=0.0063625385 laigc=-1.4681209e-011            waigc=-1.3367767e-010            paigc=4.0339002e-018 bigc=0.0018040038               wbigc=-1.4382664e-010            aigsd=0.0059804722 laigsd=-2.2470724e-011            waigsd=-1.7210843e-011            paigsd=8.5664522e-019 bigsd=0.00048472442              wbigsd=2.8664416e-011             tvoff=-0.00242207 ltvoff=1.38944e-010               wtvoff=4.06621e-010               ptvoff=-1.28635e-017 kt1=-0.69785687                lkt1=1.6794114e-008             wkt1=5.9347145e-008 pkt1=-1.8202787e-015            kt2=-0.22379967                wkt2=1.8810191e-008 ute=-2.6061728                 wute=3.237037e-007              ua1=9.9467337e-009 lua1=-3.7683439e-016            wua1=-1.3985338e-015            pua1=4.2210141e-023 ub1=-1.6474654e-17             lub1=6.2769512e-25              wub1=2.4868363e-24 pub1=-7.6747676e-32             uc1=-9.6341772e-010            luc1=3.1855103e-017 wuc1=1.4868202e-016             puc1=-4.0459477e-024            at=218841.29 lu0=-6.675631e-011             pu0=2.7836098e-018             lpdiblc2=-2.6237037e-010 wpdiblc2=-1.1005926e-009            ppdiblc2=2.9910222e-017             lbigc=-1.0689937e-011 pbigc=4.3927777e-018             lbigsd=-3.5518503e-012            pbigsd=-1.1926851e-018 lkt2=6.6080314e-009             pkt2=-7.2076676e-016            lute=7.4148148e-008 pute=-1.1964089e-014            lat=-0.0058234495              wat=-0.019008423 pat=5.5707346e-010             letab=1.3100483e-008             petab=-4.8998926e-016 leta0=5.6700699e-009             weta0=2.9845568e-009             peta0=-3.5936736e-016 lvsat=-0.0003224663              pvsat=-4.4917784e-011 jtsswgs='4.5e-007*(1+0.42*iboffp_flag_hvt)'                                jtsswgd='4.5e-007*(1+0.42*iboffp_flag_hvt)' vth0_ff=-0.0124938                 vth0_mc=0.0129012                  lvth0_ff=5.24741e-10 lvth0_mc=-5.41852e-10               wvth0_ff=1.4243e-09                 wvth0_mc=-3.56074e-09 pvth0_ff=-5.98204e-17               pvth0_mc=1.49551e-16                cit_mcl=0.00129012 lcit_mcl=-5.41852e-11               wcit_mcl=-3.56074e-10               pcit_mcl=1.49551e-17 voff_ss=0.0124938                  voff_ff=-0.011                     voff_mcl=-0.00543213 lvoff_ss=-5.24741e-10               lvoff_ff=4.62e-10                   lvoff_mcl=2.28146e-10 wvoff_ss=-1.4243e-09                wvoff_ff=-4.4e-15                   wvoff_mcl=-3.56074e-09 pvoff_ss=5.98204e-17                pvoff_ff=-3.3e-23                   pvoff_mcl=1.49551e-16 u0_ff=0.000624691                u0_mc=-0.00312346                wu0_ff=-7.12148e-11 wu0_mc=3.56074e-10                vsat_ff=-2246.91                   vsat_fs=1290.12 vsat_mcl=2580.25                    vsat_mc='9370.37-2580.25'          wvsat_ff=-0.00016185 wvsat_fs=-0.000356074               wvsat_mcl=-0.000712148               wvsat_mc='-0.00106822+0.000712148' a0_fs=-0.891358                  a0_sf=-0.950622                  la0_fs=4.33481e-08 la0_sf=3.99258e-08                wa0_fs=2.46015e-07                wa0_sf=-1.4243e-07 pa0_fs=-1.19641e-14               pa0_sf=5.98203e-15                kt1_sf=-0.0129012 lkt1_sf=5.41852e-10                wkt1_sf=3.56074e-09                pkt1_sf=-1.49551e-16 ua1_sf=-4.32716e-10               ua1_fs=7.95062e-10                ua1_ss=9.54074e-10 ua1_ff=-3.97531e-10               lua1_sf=1.31185e-17                lua1_fs=-2.6237e-17 lua1_ss=-3.14844e-17               lua1_ff=1.31185e-17                wua1_sf=5.50296e-17 wua1_fs=-9.0637e-17                wua1_ss=-1.08764e-16               wua1_ff=4.53185e-17 pua1_sf=-1.49551e-24               pua1_fs=2.99102e-24                pua1_ss=3.58923e-24 pua1_ff=-1.49551e-24               lu0_ff=-2.6237e-11                lu0_mc=1.31185e-10 pu0_ff=2.99102e-18                pu0_mc=-1.49551e-17               lvsat_ff=2.28154e-05 lvsat_fs=-5.41852e-05               lvsat_mcl=-0.00010837                lvsat_mc='-0.000393556+0.00010837' pvsat_ff=1.49551e-11                pvsat_fs=1.49551e-11                pvsat_mcl=2.99102e-11 pvsat_mc='4.48653e-11-2.99102e-11' lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_lvt_mac.global nmos ( modelid=5                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_lvt'             permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          wpemod=1 tnom=25                         toxe=1.95e-009                  toxm=1.95e-009 dtox=3.532e-010                 epsrox=3.9                        toxref=3e-009 wint=0                          lint=0                          ll=0 wl=0                          lln=1                          wln=1 lw=0                          ww=0                          lwn=1 wwn=1                          lwl=0                          wwl=0 llc=0                          wlc=0                          lwc=0 wwc=0                          lwlc=0                          wwlc=0 xl=-4e-009                    xw=6e-009                     dlc=6.25e-009 dwc=0                          dlcig=2.5e-009                   xpart=1 k1=0.292                      k3=0                          k3b=2.5 w0=0                          dvt0=1.4759776                  dvt1=1.6386118 dvt2=-0.15                      dvt0w=0                          dvt1w=0 dvt2w=0                          dsub=0.49745                    minv=-0.26054 voffl=0                          dvtp0=2.3209746e-012             dvtp1=0.1 lpe0=2.0063074e-008             lpeb=8.8958833e-009             xj=6.7e-008 ngate=2.2e+020                   ndep=1e+017                     nsd=1e+020 phin=0.13                       cdsc=0                          ud=0 cdscb=0                          cdscd=0                          nfactor=1 a1=0                          a2=1                          b0=0 b1=0                          dwg=0                          dwb=0 pdiblc1=0                          pdiblcb=1                          drout=0.56 pvag=2                          delta=0.015                      pscbe1=1e+009 pscbe2=1e-020                     fprout=300                        pdits=0 pditsd=0                          pditsl=0                          rsh=18 rdsw=86.009                     prwg=0                          prwb=0 wr=1                          alpha0=6.7554e-008                alpha1=2.7898 beta0=13.5                       agidl=5e-008                     bgidl=1.8981526e+009 cgidl=0.5                        egidl=0.31116                    bigbacc=0.0053226965 cigbacc=0.34506                    nigbacc=8.0450728                  aigbinv=0.01469171 bigbinv=0.0047951186               cigbinv=0.006                      eigbinv=1.1 nigbinv=7.0466982                  bigc=0.0011268385               cigc=-0.04 bigsd=0.00050676879              cigsd=7.6145e-020                nigc=2.7318217 poxedge=1                          pigcd=3.2220404                  ntox=1 vfbsdoff=0.01                       cgso=9.775e-011                 cgdo=9.775e-011 cgbo=0                          cgdl=1.449e-011                 cgsl=1.449e-011 clc=0                          cle=0.6                        cf='6.62e-011+9.73e-11*ccoflag_lvt' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=5                          noff=2.7                        voffcv=-0.1 tvfbsdoff=0.1                        kt1l=0                          prt=0 fnoimod=1                          tnoimod=0                          em=1.30e+007 ef=0.90                       noia=0                          noib=0 noic=0                          lintnoi=-3.79e-008                 jss=3.11e-07 jsd=3.11e-07                   jsws=9.46e-14                   jswd=9.46e-14 jswgs=9.46e-14                   jswgd=9.46e-14                   njs=1.03 njd=1.03                       ijthsfwd=0.01                       ijthdfwd=0.01 ijthsrev=0.01                       ijthdrev=0.01                       bvs=8.32 bvd=8.32                       xjbvs=1                          xjbvd=1 njtsswg=11                         xtsswgs=0.212                      xtsswgd=0.212 tnjtsswg=1                          vtsswgs=1.36                       vtsswgd=1.36 pbs=0.67                       pbd=0.67                       cjs=0.00139 cjd=0.00139                    mjs=0.313                      mjd=0.313 pbsws=0.472                      pbswd=0.472                      cjsws=1.05e-010 cjswd=1.05e-010                  mjsws=0.011                      mjswd=0.011 pbswgs=0.966                      pbswgd=0.966                      cjswgs=2.89e-010 cjswgd=2.89e-010                  mjswgs=0.643                      mjswgd=0.643 tpb=0.00113                    tcj=0.00073                    tpbsw=0.0024 tcjsw=0.00016                    tpbswg=0.00212                    tcjswg=0.00148 xtis=3                          xtid=3                          dmcg=3.8e-008 dmci=3.8e-008                   dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=2.64e-009 rshg=16.42                      gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          xrcrg1=12 xrcrg2=1                          web=2153.1                     wec=-9093.6 scref=1e-6                       kvth0we=0.00053                    k2we=0.0000 ku0we=-0.0016                    lk2we=0                          lku0we=4.5e-11 lkvth0we=-1.05e-011                 pk2we=0                          pku0we=-1e-18 pkvth0we=1.3e-018                   wk2we=0                          wku0we=3e-11 wkvth0we=-4.1e-011 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.2                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.6 bidirectionflag='bidirectionflag_mos_lvt' iboffn_flag='iboffn_flag_lvt' iboffp_flag='iboffp_flag_lvt' sigma_factor='sigma_factor_lvt' ccoflag='ccoflag_lvt' rcoflag='rcoflag_lvt' rgflag='rgflag_lvt' mismatchflag='mismatchflag_mos_lvt' globalflag='globalflag_mos_lvt' totalflag='totalflag_mos_lvt' designflag='designflag_mos_lvt' global_factor='global_factor_lvt' local_factor='local_factor_lvt' sigma_factor_flicker='sigma_factor_flicker_lvt' noiseflag='noiseflagn_lvt' noiseflag_mc='noiseflagn_lvt_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w41='2.3875*0.35355' w42='0.70711*-0.35355' w43='0.54772*0.0021707' w44='0.54772*0.81882' w45='0.54772*-0.058492' w46='0.54772*0.23016' w47='0.54772*-0.11085' w48='0.54772*-0.10416' w49='0' w50='0' tox_c='toxn_lvt'                 dxl_c='dxln_lvt'                 dxw_c='dxwn_lvt' cj_c='cjn_lvt'                  cjsw_c='cjswn_lvt'                cjswg_c='cjswgn_lvt' cgo_c='cgon_lvt'                 cgl_c='cgln_lvt'                 ddlc_c='ddlcn_lvt' ntox_c='ntoxn_lvt'                cf_c='cfn_lvt'                  dvth_c='dvthn_lvt' dlvth_c='dlvthn_lvt'               dwvth_c='dwvthn_lvt'               dpvth_c='dpvthn_lvt' du0_c='du0n_lvt'                 dlu0_c='dlu0n_lvt'                dwu0_c='dwu0n_lvt' dpu0_c='dpu0n_lvt'                dvsat_c='dvsatn_lvt'               dlvsat_c='dlvsatn_lvt' dwvsat_c='dwvsatn_lvt'              dpvsat_c='dpvsatn_lvt'              dk2_c='dk2n_lvt' dlk2_c='dlk2n_lvt'                dwk2_c='dwk2n_lvt'                dpk2_c='dpk2n_lvt' dvoff_c='dvoffn_lvt'               dlvoff_c='dlvoffn_lvt'              dwvoff_c='dwvoffn_lvt' dpvoff_c='dpvoffn_lvt'              dpdiblc2_c='dpdiblc2n_lvt'            dlpdiblc2_c='dlpdiblc2n_lvt' dwpdiblc2_c='dwpdiblc2n_lvt'           dppdiblc2_c='dppdiblc2n_lvt'           dags_c='dagsn_lvt' dlags_c='dlagsn_lvt'               dwags_c='dwagsn_lvt'               dpags_c='dpagsn_lvt' deta0_c='deta0n_lvt'               dleta0_c='dleta0n_lvt'              dweta0_c='dweta0n_lvt' dpeta0_c='dpeta0n_lvt'              dpclm_c='dpclmn_lvt'               dlpclm_c='dlpclmn_lvt' dwpclm_c='dwpclmn_lvt'              dppclm_c='dppclmn_lvt'              dminv_c='dminvn_lvt' dua1_c='dua1n_lvt'                dat_c='datn_lvt'                 dlat_c='dlatn_lvt' dwat_c='dwatn_lvt'                dpat_c='dpatn_lvt'                jtsswg_c='jtsswgn_lvt' ss_flag_c='ss_flagn_lvt'             ff_flag_c='ff_flagn_lvt'             sf_flag_c='sf_flagn_lvt' fs_flag_c='fs_flagn_lvt'             monte_flag_c='monte_flagn_lvt'         c1f_c='c1fn_lvt' c2f_c='c2fn_lvt'                 c3f_c='c3fn_lvt' global_mc='global_mc_flag_lvt' tox_g='toxn_lvt_ms_global'       dxl_g='dxln_lvt_ms_global'       dxw_g='dxwn_lvt_ms_global' cj_g='cjn_lvt_ms_global'        cjsw_g='cjswn_lvt_ms_global' cjswg_g='cjswgn_lvt_ms_global'     cgo_g='cgon_lvt_ms_global'       cgl_g='cgln_lvt_ms_global' ntox_g='ntoxn_lvt_ms_global'      cf_g='cfn_lvt_ms_global'        dvth_g='dvthn_lvt_ms_global' dlvth_g='dlvthn_lvt_ms_global'     dwvth_g='dwvthn_lvt_ms_global' dpvth_g='dpvthn_lvt_ms_global'     du0_g='du0n_lvt_ms_global'       dlu0_g='dlu0n_lvt_ms_global' dwu0_g='dwu0n_lvt_ms_global'      dpu0_g='dpu0n_lvt_ms_global' dvsat_g='dvsatn_lvt_ms_global'     dlvsat_g='dlvsatn_lvt_ms_global' dwvsat_g='dwvsatn_lvt_ms_global'    dpvsat_g='dpvsatn_lvt_ms_global' dk2_g='dk2n_lvt_ms_global'       dlk2_g='dlk2n_lvt_ms_global'      dwk2_g='dwk2n_lvt_ms_global' dpk2_g='dpk2n_lvt_ms_global'      dlvoff_g='dlvoffn_lvt_ms_global' dpvoff_g='dpvoffn_lvt_ms_global'    dpdiblc2_g='dpdiblc2n_lvt_ms_global' dags_g='dagsn_lvt_ms_global'      dwags_g='dwagsn_lvt_ms_global' dleta0_g='dleta0n_lvt_ms_global'    dpclm_g='dpclmn_lvt_ms_global' dminv_g='dminvn_lvt_ms_global'     dua1_g='dua1n_lvt_ms_global'      dat_g='datn_lvt_ms_global' ss_flag_g='ss_flagn_lvt_ms_global'   ff_flag_g='ff_flagn_lvt_ms_global' monte_flag_g='monte_flagn_lvt_ms_global'                                       sf_flag_g='sf_flagn_lvt_ms_global' fs_flag_g='fs_flagn_lvt_ms_global' weight1=-3.4493056 weight2=2.1815278 weight3=1.1797917 weight4=0.69444444 weight5=-0.48354861 tox_1=4.5194711e-012 tox_2=-9.4735394e-012 tox_3=-1.8851879e-012 tox_4=-3.747676e-011 tox_5=6.3111596e-013 dxl_1=1.0232935e-010 dxl_2=-2.1449863e-010 dxl_3=-4.2683727e-011 dxl_4=8.4852457e-010 dxl_5=1.4288909e-011 dxw_1=-6.9400556e-010 dxw_2=-8.5539453e-010 dxw_3=1.2683919e-010 dxw_4=1.8191884e-025 dxw_5=-5.8948623e-009 cj_1=9.6618e-006 cj_2=-2.1117e-006 cj_3=-2.5808e-006 cj_4=5.4672e-021 cj_5=-9.1496e-007 cjsw_1=7.2985e-013 cjsw_2=-1.5952e-013 cjsw_3=-1.9495e-013 cjsw_4=4.1299e-028 cjsw_5=-6.9116e-014 cjswg_1=2.0088e-012 cjswg_2=-4.3905e-013 cjswg_3=-5.3658e-013 cjswg_4=1.1367e-027 cjswg_5=-1.9023e-013 cgo_1=-6.7946e-013 cgo_2=1.485e-013 cgo_3=1.8149e-013 cgo_4=-7.277e-028 cgo_5=6.4344e-014 cgl_1=-1.0072e-013 cgl_2=2.2013e-014 cgl_3=2.6903e-014 cgl_4=1.6431e-029 cgl_5=9.538e-015 ntox_1=-0.0017541 ntox_2=0.00053405 ntox_3=-0.0086448 ntox_4=2.8165e-018 ntox_5=-4.685e-005 cf_1=-4.6015e-013 cf_2=1.0057e-013 cf_3=1.2291e-013 cf_4=-8.8346e-029 cf_5=4.3576e-014 dvth_1=0.0033089 dvth_2=0.0042337 dvth_3=-0.00067301 dvth_4=-7.3914e-018 dvth_5=-0.00090171 dlvth_1=5.8065e-011 dlvth_2=8.3376e-011 dlvth_3=-7.8345e-012 dlvth_4=1.5904e-025 dlvth_5=-1.7489e-011 dwvth_1=2.3254e-010 dwvth_2=1.2765e-010 dwvth_3=-9.9243e-011 dwvth_4=-1.6633e-025 dwvth_5=-4.5047e-011 dpvth_1=1.307e-017 dpvth_2=9.2039e-018 dpvth_3=5.3295e-019 dpvth_4=3.0253e-033 dpvth_5=-2.4723e-018 du0_1=0.0001025 du0_2=0.00028777 du0_3=-1.9725e-005 du0_4=-5.5691e-020 du0_5=-5.4776e-005 dlu0_1=5.329e-013 dlu0_2=6.5617e-012 dlu0_3=3.8759e-013 dlu0_4=6.5199e-027 dlu0_5=-1.0039e-012 dwu0_1=7.8655e-012 dwu0_2=3.9425e-011 dwu0_3=-3.4395e-012 dwu0_4=-2.3814e-026 dwu0_5=-6.8346e-012 dpu0_1=5.8454e-020 dpu0_2=1.516e-018 dpu0_3=1.8e-019 dpu0_4=6.8821e-034 dpu0_5=-2.8381e-019 dvsat_1=184.3 dvsat_2=2148.3 dvsat_3=-63.191 dvsat_4=6.7623e-013 dvsat_5=-380.24 dlvsat_1=5.6747e-005 dlvsat_2=-1.2768e-005 dlvsat_3=6.9746e-006 dlvsat_4=9.8966e-022 dlvsat_5=-4.8567e-006 dwvsat_1=5.4084e-005 dwvsat_2=0.00063946 dwvsat_3=-3.7941e-005 dwvsat_4=-1.7722e-019 dwvsat_5=-0.00012226 dpvsat_1=-2.7789e-012 dpvsat_2=6.9129e-013 dpvsat_3=-4.3352e-012 dpvsat_4=-1.0447e-027 dpvsat_5=1.445e-013 dk2_1=0.00031302 dk2_2=-7.7023e-005 dk2_3=0.00043715 dk2_4=-4.6222e-019 dk2_5=-1.7473e-005 dlk2_1=5.846e-012 dlk2_2=-1.5532e-012 dlk2_3=1.5103e-011 dlk2_4=3.9401e-027 dlk2_5=-1.642e-013 dwk2_1=3.2416e-011 dwk2_2=-7.5906e-012 dwk2_3=2.1936e-011 dwk2_4=7.1397e-027 dwk2_5=-2.3548e-012 dpk2_1=2.5768e-018 dpk2_2=-5.8299e-019 dpk2_3=5.0945e-019 dpk2_4=-1.902e-033 dpk2_5=-2.1603e-019 dlvoff_1=-1.7188e-011 dlvoff_2=3.649e-012 dlvoff_3=1.1101e-011 dlvoff_4=3.9191e-028 dlvoff_5=1.7798e-012 dpvoff_1=6.2655e-018 dpvoff_2=-1.2617e-018 dpvoff_3=-8.1831e-018 dpvoff_4=1.3985e-034 dpvoff_5=-7.4545e-019 dpdiblc2_1=-7.7454e-005 dpdiblc2_2=1.6928e-005 dpdiblc2_3=2.0689e-005 dpdiblc2_4=2.8334e-020 dpdiblc2_5=7.3348e-006 dags_1=0.050814 dags_2=0.034103 dags_3=-0.0047103 dags_4=-4.0574e-017 dags_5=-0.0091442 dwags_1=1.0031e-009 dwags_2=-4.7467e-009 dwags_3=-1.9162e-009 dwags_4=7.6751e-024 dwags_5=3.9134e-010 dleta0_1=-1.986e-011 dleta0_2=4.3405e-012 dleta0_3=5.3048e-012 dleta0_4=-9.2964e-027 dleta0_5=1.8807e-012 dpclm_1=-0.00993 dpclm_2=0.0021703 dpclm_3=0.0026524 dpclm_4=-1.6229e-017 dpclm_5=0.00094035 dminv_1=-0.004965 dminv_2=0.0010851 dminv_3=0.0013262 dminv_4=-3.516e-018 dminv_5=0.00047018 dua1_1=3.972e-012 dua1_2=-8.6811e-013 dua1_3=-1.061e-012 dua1_4=-5.7089e-027 dua1_5=-3.7614e-013 dat_1=1489.5 dat_2=-325.54 dat_3=-397.86 dat_4=-8.3233e-013 dat_5=-141.05 ss_flag_1=0.05343 ss_flag_2=-0.01383 ss_flag_3=0.11592 ss_flag_4=-7.8776e-018 ss_flag_5=-0.0020174 ff_flag_1=-0.04587 ff_flag_2=0.0078727 ff_flag_3=0.14244 ff_flag_4=-6.1309e-017 ff_flag_5=0.0073861 monte_flag_1=0.085275 monte_flag_2=-0.17875 monte_flag_3=-0.03557 monte_flag_4=0.707108 monte_flag_5=0.0119075 sigma_local=1                          a_1=0.955086 b_1=-0.00272346                c_1=-0.000561476               d_1=0.000343593 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1.06037                    b_2=-0.00133227                c_2=-0.00624525 d_2=-0.00057247                a_3=1.01463                    b_3=-0.00527586 c_3=-0.0081346                 d_3=-0.00020372                e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.8 b_4=0.0002                     c_4=-0.0075                    d_4=-0.00003 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=0.74                       b_5=-2.5e-3                    c_5=-0.0075 d_5=-0.00003                   e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.0026                     mis_a_2=0.08                       mis_a_3=0.07 mis_b_1=0.0033                     mis_b_2=0.08                       mis_b_3=0.00 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.00080                    mis_d_2=0.00                       mis_d_3=0 mis_e_1=0.0024                     mis_e_2=-0.09                      mis_e_3=0 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-4e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18 cf0=6.62e-011                  cco=9.73e-11 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.4                        l_rjtsswg=3e-5                       ll_rjtsswg=3 w_rjtsswg=0                          ww_rjtsswg=0                          p_rjtsswg=0.0 noimod=1                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6                sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=0                   lreflod=1e-6                llodref=3 lod_clamp=-1e90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=1 kvth00=0                   lkvth00=0                   wkvth00=0 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0 lodeta00=1 wlod00=0 ku000=0                   lku000=0                   wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0                   lkvth000=0                   wkvth000=0         		pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=0                   wku01=0 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=0                   wkvth01=0 pkvth01=0                   llodvth1=1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.06               lku02=1.5e-7              wku02=7e-8 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=-0.5 kvth02=7e-3                lkvth02=-9e-9               wkvth02=16e-9 pkvth02=1e-15               llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=-0.03               lku03=7e5                 wku03=-5e-8 pku03=0                   tku03=0                   llodku03=-1 wlodku03=1                   kvsat3=0 kvth03=9e-3                lkvth03=-3e-9               wkvth03=-2e-8 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=-0.000                   lku003=-0.0e-9                   wku003=-0e-9         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0.0e-3                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl='0.15*01'           wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl='1.4e-12*1'         ldplkvth0=1.5                 pkvth0dpl=0.0e-19 ku0dpl='0.50*0'            wku0dpl=0e-8                wdplku0=1 lku0dpl=5.0e-8              ldplku0=1.0                 pku0dpl=0.0e-11 keta0dpl='0.07*0'            wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0.00                wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.000              wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx='0.25*1'            wku0dpx=0e-9                wdpxku0=1 lku0dpx='1.0e-8*1'          ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps='0.1*1'             wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='-0.70*1'           wku0dps=-0.0e-9             wdpsku0=1 lku0dps='9.0e-15*1'         ldpsku0=2.0                 pku0dps='-7.0e-23*0' keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps='-0.3*0'            wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa='0.01*0'            wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa='1.0e-9*0'          ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa='0.050*0'           wku0dpa=0e-7                wdpaku0=1 lku0dpa=0.0e-11             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=-0.0                wka0dpa=0                   wdpaka0=1 lka0dpa=-0.0e-7             ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa='1.5*0'             wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2='0.005*1'           wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2='3e-9*1'            ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.000               wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2='2.5e-5*1'          ldp2ku0=0.5                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2='0.5*0'             wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx='0.050*2'           wkvth0enx='8.0e-9*1'          wenxkvth0=1 lkvth0enx='1.0e-8*1'          lenxkvth0=1.0                 pkvth0enx=0 ku0enx='-0.90*1.7'         wku0enx='-0.9e-8*1.5'       wenxku0=1 lku0enx='2.0e-7*1'          lenxku0=1.0                 pku0enx='-3.0e-16*1.7' keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0.0                 wka0enx=0                   wenxka0=1 lka0enx='1.0e-7*2'          lenxka0=1.0                 pka0enx='1.0e-14*1.7' kvsatenx=-0.0                wenx=0                   ku0enx0='0.15*0' eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.01e-6 kvth0eny='0.04*1.7'          wkvth0eny='4.0e-10*4'         wenykvth0=1 lkvth0eny='1.0e-7*1.7'        lenykvth0=1.0                 pkvth0eny=0 ku0eny='-0.70*2'           wku0eny='-1.1e-8*1'         wenyku0=1 ku0eny0='0.025*0'           wku0eny0=0                   weny0ku0=1 lku0eny='6.0e-10*1.7'       lenyku0=1.5                 pku0eny=-0.0e-14 keta0eny=0.00                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-8             wenyka0=1 lka0eny='-6.0e-8*1.7'       lenyka0=1.0                 pka0eny='1.0e-14*1.7' kvsateny=-0.0                weny=0 kvth0eny1=0.000              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=0 ku0eny1='0.15*1.7'         wku0eny1=0.0e-8             weny1ku0=1 lku0eny1='1.0e-5*1.4'       leny1ku0=1.0                pku0eny1=-0.0e-14 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1.0                pka0eny1=0 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=-0.045              wkvth0rx=-0.0e-5             wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0.0e-16 ku0rx='0.3'               wku0rx=0.0e-8              wrxku0=1.0 lku0rx='-3.5e-10*0'        lrxku0=1                   pku0rx=0.0e-15 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.0                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=0.9027e-5           ringymin=0.117e-6 kvth0ry='-0.03*1'           wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry=0.0e-8              lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry='-0.02*1'           wku0ry=-0.0e-8             wryku0=1.0 lku0ry='-1.0e-8*1'         lryku0=1.0                 pku0ry=-0.0e-16 keta0ry=0.00                wketa0ry=0                   wryketa0=1 kvsatry=0                   wry=0 kvth0ry0=0.01                ku0ry0=0.02 sfxref=9.0e-8            sfxmax=3.906e-6           minwodx=0.0e-6 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0009            lkvth0odx1b=0.0e-7            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.0028           lku0odx1b=0.8e-10           lodx1bku0=1.0 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6              sfymax=10e-6             minwody=0.9e-6 wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-1.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.000            lkvth0odyb=0.0e-10           lodybkvth0=1.0 wkvth0odyb=-2.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.03             lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-1.0e-7           wodybku0=1.0               pku0odyb=0 web_mac=0  wec_mac=0 kvsatwe=0.0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model nch_lvt_mac.1 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=9.01e-06                   vth0=0.35295609 lvth0=3.3798175e-008             wvth0=-1.2642487e-008            pvth0=-1.3753726e-014 k2=0.012533395                lk2=2.6446003e-013             wk2=-1.1531474e-008 pk2=-2.3981175e-019            cit=0.0024549256               lcit=-3.9648754e-010 wcit=3.70639e-010               pcit=-1.6256474e-016            voff=-0.1384174 lvoff=-2.9025039e-008            wvoff=-1.2719601e-008            pvoff=7.2630841e-015 eta0=0.0072237037               weta0=-2.0146756e-009            etab=-0.03571197 wetab=-1.8938152e-010            u0=0.018406123                wu0=6.5498009e-010 ua=-1.4758974e-009            lua=-1.1180314e-017            wua=3.2643736e-017 pua=-2.9930087e-023            ub=1.8755037e-018             lub=-8.2631857e-027 wub=-1.1798396e-027            pub=7.4864462e-033             uc=1.3842061e-010 wuc=-3.3605393e-017            vsat=120000                     a0=3.3059527 la0=-5.5871247e-007            wa0=-4.2565447e-007            pa0=2.7687944e-013 ags=1.2275722                  lags=6.5320872e-007             wags=2.8873715e-008 pags=-1.5092742e-013            keta=-0.077926708               lketa=-6.37287e-008 wketa=4.2356802e-008             pketa=2.492496e-014              pclm=0.26792894 lpclm=1.8788935e-007             wpclm=8.9590604e-008             ppclm=1.0024399e-013 pdiblc2=0.0014023181               lpdiblc2=8.7874663e-010             wpdiblc2=1.301521e-011 ppdiblc2=-1.1708483e-016            aigbacc=0.013336995                laigbacc=8.9264994e-011 waigbacc=1.6627931e-011             paigbacc=-2.7816816e-017            aigc=0.010776112 laigc=-9.6981495e-011            waigc=4.4778023e-011             paigc=4.6531202e-017 aigsd=0.0097031278               laigsd=6.6969716e-011             waigsd=2.5737952e-011 paigsd=3.588756e-018              tvoff=0.00194164                 ltvoff=-1.73382e-010 wtvoff=-2.04096e-010              ptvoff=2.36432e-017               kt1=-0.17475901 lkt1=-1.1011332e-012            wkt1=1.0707816e-008             pkt1=2.8368345e-018 kt2=-0.059088294               lkt2=-9.9511311e-016            wkt2=-8.2099056e-009 pkt2=1.8956347e-029             ute=-1.2070146                 lute=-1.1064183e-013 wute=2.2435698e-007             pute=1.002415e-019              ua1=1.3753943e-009 lua1=1.4085568e-016             wua1=9.6075649e-017             pua1=-1.3933569e-022 ub1=-1.164586e-018             lub1=-2.492314e-025             wub1=2.6396124e-025 pub1=1.1185774e-031             uc1=6.9675516e-011             luc1=-6.5684066e-017 wuc1=9.4694261e-017             puc1=9.021706e-024              at=140000 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' lu0=0                          pu0=0                          lat=0 wat=0                          pat=0                          lvsat=0 wvsat=0                          pvsat=0                          leta0=0 peta0=0                          a0_fs=0.00122973                 la0_fs=-1.10639e-08 wa0_fs=-1.11414e-09               pa0_fs=1.00239e-14                ags_ff=0.259165 ags_fs=0.203635                   ags_ss=-0.271586                  ags_sf=-0.209845 lags_ff=-2.32212e-07               lags_fs=-1.82456e-07               lags_ss=2.43341e-07 lags_sf=1.88021e-07                wags_ff=-3.35622e-08               wags_fs=-3.35621e-08 wags_ss=1.45436e-07                wags_sf=8.94991e-08                pags_ff=3.0072e-14 pags_fs=3.00715e-14                pags_ss=-1.30311e-13               pags_sf=-8.0191e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.2 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.38522647 lvth0=4.8839139e-009             wvth0=-3.6149052e-008            pvth0=7.308156e-015 k2=0.018946718                lk2=-5.746073e-009             wk2=-1.2470335e-008 pk2=8.4098043e-016             cit=0.0019979873               lcit=1.2929162e-011 wcit=4.8023987e-010             pcit=-2.6076712e-016            voff=-0.17059922 lvoff=-1.9012832e-010            wvoff=-1.7093867e-009            pvoff=-2.6020677e-015 eta0=0.0072237037               weta0=-2.0146756e-009            etab=-0.035711993 wetab=-1.8917086e-010            u0=0.018346924                wu0=6.9375931e-010 ua=-1.4506328e-009            lua=-3.3817438e-017            wua=-2.7693963e-018 pua=1.8000797e-024             ub=1.9065332e-018             lub=-3.6065608e-026 wub=2.0073588e-026             pub=-1.1556625e-032            uc=1.3366189e-010 wuc=-1.9630155e-017            vsat=120000                     a0=2.6989741 la0=-1.4859698e-008            wa0=2.9122618e-007             pa0=-3.6544562e-013 ags=1.3105252                  lags=5.7888287e-007             wags=-1.0718441e-007 pags=-2.901934e-014             keta=-0.16828175                lketa=1.7229415e-008 wketa=9.806299e-008              pketa=-2.4987784e-014            pclm=0.42114975 lpclm=5.0603503e-008             wpclm=2.5263833e-007             ppclm=-4.5846773e-014 pdiblc2=0.002145881                lpdiblc2=2.1251428e-010             wpdiblc2=-3.4597047e-011 ppdiblc2=-7.4424247e-017            aigbacc=0.013249633                laigbacc=1.6754167e-010 waigbacc=-1.1364965e-011            paigbacc=-2.7351815e-018            aigc=0.010677784 laigc=-8.8788269e-012            waigc=1.4479622e-010             paigc=-4.3085102e-017 aigsd=0.0098121141               laigsd=-3.0682053e-011            waigsd=4.5575857e-011 paigsd=-1.4186008e-017            tvoff=0.00194352                 ltvoff=-1.75061e-010 wtvoff=-3.81489e-010              ptvoff=1.82588e-016               kt1=-0.1756879 lkt1=8.3118978e-010             wkt1=1.9776312e-009             pkt1=7.8250826e-015 kt2=-0.055987658               lkt2=-2.7781706e-009            wkt2=-1.3988334e-008 pkt2=5.1774715e-015             ute=-1.1910526                 lute=-1.4302097e-008 wute=2.5179527e-007             pute=-2.4584608e-014            ua1=1.9129953e-009 lua1=-3.4083482e-016            wua1=-1.5983021e-016            pua1=8.9955964e-023 ub1=-1.7533599e-018            lub1=2.7831005e-025             wub1=7.7924276e-025 pub1=-3.498345e-031             uc1=-2.3924675e-011            luc1=1.8181706e-017 wuc1=1.4469847e-016             puc1=-3.578207e-023             at=140554.29 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=2.0958297e-014             petab=-1.8875042e-019            lu0=5.3041964e-011 pu0=-3.474618e-017             luc=4.2638112e-018             puc=-1.2521813e-023 lat=-0.00049664211             wat=-0.0049919183              pat=4.4727588e-009 lvsat=0                          wvsat=0                          pvsat=0 leta0=0                          peta0=0                          a0_ff=-0.495556 a0_ss=0.495556                   a0_fs=-0.154178                  a0_sf=0.330262 la0_ff=4.44018e-07                la0_ss=-4.44018e-07               la0_fs=1.28181e-07 la0_sf=-2.95915e-07               wa0_ff=3.7e-13                    wa0_ss=-3.7e-13 wa0_fs=-1.29698e-07               wa0_sf=1.49756e-07                pa0_ff=3.3e-19 pa0_ss=-3.3e-19                   pa0_fs=1.25235e-13                pa0_sf=-1.34181e-13 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.3 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.39936644 lvth0=-1.4225107e-009            wvth0=-1.7099367e-008            pvth0=-1.1880033e-015 k2=0.012911792                lk2=-3.0544961e-009            wk2=-9.4670502e-009 pk2=-4.984848e-016             cit=0.0021333744               lcit=-4.7453457e-011 wcit=-6.7810164e-010            pcit=2.558532e-016              voff=-0.16599878 lvoff=-2.241924e-009             wvoff=-8.5992483e-009            pvoff=4.7081058e-016 eta0=0.0072237037               weta0=-2.0146756e-009            etab=-0.036126381 wetab=3.5338374e-009             u0=0.018343162                wu0=5.5864755e-010 ua=-1.4504207e-009            lua=-3.3912024e-017            wua=1.9628807e-017 pua=-8.1895189e-024            ub=1.8277213e-018             lub=-9.1550252e-028 wub=1.0224139e-026             pub=-7.1637705e-033            uc=1.5403533e-010 wuc=-4.2550466e-017            vsat=120000                     a0=3.5922807 la0=-4.1327442e-007            wa0=-9.5094971e-007            pa0=1.8856483e-013 ags=1.684636                   lags=4.1202947e-007             wags=7.1747913e-007 pags=-3.9681928e-013            keta=-0.12248874                lketa=-3.1942661e-009 wketa=3.7048159e-008             pketa=2.2248304e-015             pclm=0.36544889 lpclm=7.5446084e-008             wpclm=2.0131133e-007             ppclm=-2.2954933e-014 pdiblc2=0.0025388149               lpdiblc2=3.726573e-011              wpdiblc2=-2.648954e-010 ppdiblc2=2.8288817e-017             aigbacc=0.013677124                laigbacc=-2.3119205e-011 waigbacc=-1.8886682e-010            paigbacc=7.6430645e-017             aigc=0.010664967 laigc=-3.1628224e-012            waigc=3.9994051e-011             paigc=3.6566654e-018 aigsd=0.0097098084               laigsd=1.4946316e-011             waigsd=1.2134043e-011 paigsd=7.2904149e-019             tvoff=0.00163525                 ltvoff=-3.7573e-011 wtvoff=1.16963e-010               ptvoff=-3.97218e-017              kt1=-0.18394877 lkt1=4.515536e-009              wkt1=3.4789394e-008             pkt1=-6.8089636e-015 kt2=-0.055667846               lkt2=-2.9208068e-009            wkt2=-2.0492051e-009 pkt2=-1.4737985e-016            ute=-1.2368404                 lute=6.1192452e-009 wute=3.5336926e-007             pute=-6.9886607e-014            ua1=1.6833409e-009 lua1=-2.3840897e-016            wua1=4.9103293e-018             pua1=1.6481684e-023 ub1=-1.7773779e-018            lub1=2.8902209e-025             wub1=2.1570983e-025 pub1=-9.849882e-032             uc1=-6.2122646e-011            luc1=3.5218001e-017 wuc1=1.2287799e-016             puc1=-2.6050134e-023            at=190696.58 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=1.8483786e-010             petab=-1.6606504e-015            lu0=5.4719708e-011 pu0=2.5513664e-017             luc=-4.822743e-018             puc=-2.2993541e-024 lat=-0.022860106               wat=0.01441469                 pat=-4.1825883e-009 lvsat=0                          wvsat=0                          pvsat=0 leta0=0                          peta0=0                          vsat_ff=3775.92 vsat_ss=-2717.95                   vsat_fs=1811.96                    vsat_sf=-1811.96 a0_ff=0.308669                   a0_ss=-0.499998                  a0_fs=-0.0178713 a0_sf=-0.453924                  la0_ff=8.53329e-08                la0_ss=-2.91e-13 la0_fs=6.73888e-08                la0_sf=5.38322e-08                wa0_ff=9.12623e-08 wa0_ss=-2.6e-13                   wa0_fs=2.87991e-07                wa0_sf=-2.87991e-07 pa0_ff=-4.0703e-14                pa0_ss=-1.4e-19                   pa0_fs=-6.10545e-14 pa0_sf=6.10543e-14                lvsat_ff=-0.00168405                lvsat_ss=0.00121221 lvsat_fs=-0.000808137               lvsat_sf=0.000808137                wvsat_ff=-0.00136893 wvsat_ss=1.6e-09                    wvsat_fs=-1.1e-09                   wvsat_sf=1.1e-09 pvsat_ff=6.10539e-10                pvsat_ss=4.9e-15                    pvsat_fs=4.3e-16 pvsat_sf=-4.3e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.4 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.40952708 lvth0=-3.5765667e-009            wvth0=-3.0359966e-008            pvth0=1.6232436e-015 k2=-0.0087843714              lk2=1.5450906e-009             wk2=-4.9857823e-009 pk2=-1.4485136e-015            cit=0.00050265364              lcit=2.9825934e-010 wcit=1.2515839e-009             pcit=-1.5324013e-016            voff=-0.17256781 lvoff=-8.492903e-010             wvoff=-1.9220586e-009            pvoff=-9.4475363e-016 eta0=0.0072237037               weta0=-2.0146756e-009            etab=-0.014224829 wetab=-1.6215057e-008            u0=0.018632629                wu0=7.4049e-010 ua=-1.6585866e-009            lua=1.021914e-017              wua=-4.8932047e-017 pua=6.3453822e-024             ub=1.8474791e-018             lub=-5.1041387e-027 wub=2.9222093e-026             pub=-1.1191337e-032            uc=1.1161013e-010 wuc=-3.6041708e-017            vsat=123148.63                  a0=3.7960492 la0=-4.5647333e-007            wa0=5.0531507e-007             pa0=-1.2016331e-013 ags=4.056923                   lags=-9.0895376e-008            wags=-1.9421722e-006 pags=1.670268e-013              keta=-0.11440005                lketa=-4.909068e-009 wketa=7.2891985e-008             pketa=-5.3740606e-015            pclm=0.3652947 lpclm=7.5478773e-008             wpclm=1.0524059e-007             ppclm=-2.587937e-015 pdiblc2=0.0028070477               lpdiblc2=-1.9599619e-011            wpdiblc2=1.3273544e-011 ppdiblc2=-3.0682998e-017            aigbacc=0.013945844                laigbacc=-8.0087949e-011 waigbacc=5.5941312e-011             paigbacc=2.4531321e-017             aigc=0.010624409 laigc=5.4356444e-012             waigc=1.013022e-010              paigc=-9.340662e-018 aigsd=0.009857962                laigsd=-1.6462255e-011            waigsd=2.3028984e-011 paigsd=-1.580686e-018             tvoff=0.00157197                 ltvoff=-2.41571e-011 wtvoff=-3.62955e-010              ptvoff=6.20208e-017               kt1=-0.16007341 lkt1=-5.460398e-010             wkt1=-1.6753838e-008            pkt1=4.1182016e-015 kt2=-0.068963192               lkt2=-1.0219339e-010            wkt2=-5.5486326e-009 pkt2=5.9449877e-016             ute=-1.2083324                 lute=7.5563773e-011 wute=1.7624532e-008             pute=1.2912748e-015             ua1=7.1787326e-010 lua1=-3.3729831e-017            wua1=2.4151349e-016             pua1=-3.3678186e-023 ub1=-2.8723079e-019            lub1=-2.6889101e-026            wub1=-6.0749112e-025 pub1=7.6019782e-032             uc1=1.301165e-010              luc1=-5.5366972e-018 wuc1=-3.8502688e-017            puc1=8.1625699e-024             at=84503.669 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-4.458291e-009             petab=2.5261151e-015             lu0=-6.6471352e-012 pu0=-1.3036936e-017            luc=4.1713981e-018             puc=-3.6792109e-024 lat=-0.00034720806             wat=0.0080428192               pat=-2.8317518e-009 lvsat=-0.00066751032             wvsat=0.0020763524               pvsat=-4.401867e-010 leta0=0                          peta0=0                          vsat_ff=-7012.42 vsat_ss=5123.94                    vsat_fs=-3365.08                   vsat_sf=3365.08 a0_ff=1.12834                    a0_ss=-0.765383                  a0_fs=0.466817 a0_sf=-0.260621                  la0_ff=-8.84375e-08               la0_ss=5.62611e-08 la0_fs=-3.53655e-08               la0_sf=1.28515e-08                wa0_ff=-1.69495e-07 wa0_ss=-6.87544e-08               wa0_fs=3.43774e-08                wa0_sf=-6.8754e-08 pa0_ff=1.4576e-14                 pa0_ss=1.45758e-14                pa0_fs=-7.28791e-15 pa0_sf=1.45758e-14                lvsat_ff=0.000603068                lvsat_ss=-0.000450279 lvsat_fs=0.000289396                lvsat_sf=-0.000289396               wvsat_ff=0.0025423 wvsat_ss=-0.000687535               wvsat_fs=5e-10                      wvsat_sf=-5e-10 pvsat_ff=-2.18637e-10               pvsat_ss=1.45758e-10                pvsat_fs=-2.7e-16 pvsat_sf=2.7e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.5 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.37412592 lvth0=-5.3206665e-010            wvth0=-2.1932243e-008            pvth0=8.9845951e-016 k2=0.0091911182               lk2=-8.0151897e-013            wk2=-2.4428151e-008 pk2=2.2353017e-016             cit=0.0022947729               lcit=1.4413708e-010 wcit=-8.0672312e-010            pcit=2.3774268e-017             voff=-0.16461842 lvoff=-1.5329376e-009            wvoff=-1.5172889e-008            pvoff=1.9481783e-016 eta0=0.0008079103               weta0=-1.1599299e-008            etab=-0.10629476 wetab=1.4333139e-008             u0=0.019784759                wu0=2.1748809e-010 ua=-1.7065146e-009            lua=1.4340946e-017             wua=9.9431609e-018 pua=1.2821143e-024             ub=1.7213377e-018             lub=5.744021e-027 wub=8.4769959e-027             pub=-9.4072584e-033            uc=7.7652678e-011 wuc=-2.2844882e-017            vsat=97695.04                   a0=2.1690967 la0=-3.1655542e-007            wa0=-2.5827556e-006            pa0=1.4541076e-013 ags=3                          lags=-1.3360083e-015            wags=-2.406418e-013 pags=1.203209e-020              keta=-0.24513912                lketa=6.3344916e-009 wketa=4.424824e-008              pketa=-2.9106986e-015            pclm=1.5803922 lpclm=-2.9019612e-008            wpclm=1.7952095e-007             ppclm=-8.9760475e-015 pdiblc2=0.0026113941               lpdiblc2=-2.7734074e-012            wpdiblc2=-1.2105636e-010 ppdiblc2=-1.9130626e-017            aigbacc=0.013110116                laigbacc=-8.2152869e-012 waigbacc=5.8525501e-010             paigbacc=-2.0989656e-017            aigc=0.010742555 laigc=-4.724926e-012             waigc=-1.2413591e-012            paigc=-5.2191597e-019 aigsd=0.0096677679               laigsd=-1.0556545e-013            waigsd=-1.3035986e-012 paigsd=5.119161e-019              tvoff=0.000796787                ltvoff=4.25082e-011 wtvoff=1.04629e-009               ptvoff=-5.91746e-017              kt1=-0.20817554 lkt1=3.5907435e-009             wkt1=4.7028222e-008             pkt1=-1.3670555e-015 kt2=-0.084044333               lkt2=1.1947847e-009             wkt2=1.3997659e-009 pkt2=-3.0634905e-018            ute=-1.4693145                 lute=2.2520022e-008 wute=1.1509271e-008             pute=1.8171873e-015             ua1=-2.4905519e-010 lua1=4.9426016e-017             wua1=3.8318733e-016             pua1=-4.5862137e-023 ub1=-3.9847015e-019            lub1=-1.7322515e-026            wub1=3.2282919e-026 pub1=2.0999215e-032             uc1=2.9917366e-011             luc1=3.080428e-018 wuc1=7.8796199e-017             puc1=-1.9251344e-024            at=118766.67 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=3.459723e-009              petab=-1.0102973e-016            lu0=-1.0573031e-010 pu0=3.1941229e-017             luc=7.0917392e-018             puc=-4.8141379e-024 lat=-0.0032938259              wat=-0.080976266               pat=4.8238896e-009 lvsat=0.0015214987               wvsat=-0.012927586               pvsat=8.5015199e-010 leta0=5.5175823e-010             peta0=8.2427763e-016             vsat_ss=2821.27 vsat_ff=-310.661                   a0_ff=0.238889                   a0_ss=-0.265606 a0_fs=0.132803                   a0_sf=-0.265606                  la0_ff=-1.19445e-08 la0_ss=1.32803e-08                la0_fs=-6.64014e-09               la0_sf=1.32803e-08 wa0_ff=-1.9e-13                   wa0_ss=2.40639e-07                wa0_fs=-1.20319e-07 wa0_sf=2.40639e-07                pa0_ff=-4.1e-20                   pa0_ss=-1.20319e-14 pa0_fs=6.01597e-15                pa0_sf=-1.20319e-14               lvsat_ss=-0.000252248 lvsat_ff=2.67169e-05                wvsat_ss=-0.000391742               wvsat_ff=0.00279813 pvsat_ss=1.2032e-10                 pvsat_ff=-2.40639e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.6 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.35373028 lvth0=4.8771522e-010             wvth0=5.3551893e-009             pvth0=-4.6591212e-016 k2=-0.01470946                lk2=1.1942274e-009             wk2=-1.7938561e-008 pk2=-1.0094934e-016            cit=-0.0027865798              lcit=3.9820471e-010 wcit=3.318169e-009              pcit=-1.8247034e-016            voff=-0.11892108 lvoff=-3.8178049e-009            wvoff=-5.4796394e-008            pvoff=2.175993e-015 eta0=-0.015122861               weta0=1.7398852e-008             etab=-0.089885756 wetab=5.2390517e-008             u0=0.019342574                wu0=5.5743218e-010 ua=-1.5122627e-009            lua=4.6283537e-018             wua=-3.0271398e-016 pua=1.6914972e-023             ub=1.7552851e-018             lub=4.0466505e-027 wub=7.8361039e-026             pub=-1.2901461e-032            uc=1.1070311e-010 wuc=-1.39324e-016              vsat=71394.118                  a0=-4.1200472 la0=-2.0982281e-009            wa0=1.3573368e-005             pa0=-6.6239542e-013 ags=3                          lags=0                          wags=0 pags=0                          keta=-0.16752094                lketa=2.4535827e-009 wketa=1.7700254e-008             pketa=-1.5832992e-015            pclm=1.4555551 lpclm=-2.277776e-008             wpclm=0                          ppclm=0 pdiblc2=0.0025559259               lpdiblc2=0                          wpdiblc2=-5.0366889e-010 ppdiblc2=0                          aigbacc=0.01459125                 laigbacc=-8.2272002e-011 waigbacc=2.3326961e-010             paigbacc=-3.3903867e-018            aigc=0.010840735 laigc=-9.6339374e-012            waigc=-9.141512e-012             paigc=-1.2690833e-019 aigsd=0.0093811246               laigsd=1.4226601e-011             waigsd=-6.5424484e-012 paigsd=7.7385859e-019             tvoff=0.00342212                 ltvoff=-8.87585e-011 wtvoff=-1.95053e-010              ptvoff=2.89271e-018               kt1=-0.070576438 lkt1=-3.2892118e-009            wkt1=6.3705418e-008             pkt1=-2.2009154e-015 kt2=-0.062497294               lkt2=1.1743276e-010             wkt2=2.2488147e-008 pkt2=-1.0574825e-015            ute=-1.5472144                 lute=2.6415016e-008 wute=5.5523528e-007             pute=-2.5369113e-014            ua1=9.7594558e-010 lua1=-1.1824023e-017            wua1=-2.3579667e-015            pua1=9.1195565e-023 ub1=-2.4891723e-018            lub1=8.7212591e-026             wub1=4.4092278e-024 pub1=-1.9784803e-031            uc1=-2.4486979e-010            luc1=1.6819786e-017 wuc1=4.4412403e-016             puc1=-2.0191526e-023            at=-62342.206 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=2.6392728e-009             petab=-2.0038986e-015            lu0=-8.3621074e-011 pu0=1.4944024e-017             luc=5.4392174e-018             puc=1.0098179e-024 lat=0.0057616177               wat=0.095138039                pat=-3.9818257e-009 lvsat=0.0028365448               wvsat=0.047767415                pvsat=-2.1845981e-009 leta0=1.3482968e-009             peta0=-6.2562994e-016            vsat_ff=10353.7 vsat_ss=-32614                     vsat_fs=5065.04                    lvsat_ff=-0.000506504 lvsat_ss=0.00151951                 lvsat_fs=-0.000253252               wvsat_ff=-0.0111925 wvsat_ss=0.0295483                  wvsat_fs=-0.00458893                pvsat_ff=4.58893e-10 pvsat_ss=-1.37668e-09               pvsat_fs=2.29446e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.7 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=9e-007                     wmax=9.01e-06                   vth0=0.39327703 lvth0=-1.1337015e-009            wvth0=-1.6054095e-008            pvth0=4.1186851e-016 k2=0.055831994                lk2=-1.6979722e-009            wk2=-3.4697125e-008 pk2=5.8615177e-016             cit=0.001902246                lcit=2.0596285e-010 wcit=-5.7675801e-009            pcit=1.9004537e-016             voff=-0.12216855 lvoff=-3.6846584e-009            wvoff=-1.4876312e-008            pvoff=5.392697e-016 eta0=-0.014099892               weta0=1.6910291e-008             etab=-0.045860636 wetab=3.3617755e-009             u0=0.018431765                wu0=1.2381619e-009 ua=-1.6044085e-009            lua=8.4063308e-018             wua=-1.1399636e-017 pua=4.9710832e-024             ub=1.6900104e-018             lub=6.7229121e-027 wub=6.8373537e-026             pub=-1.2491973e-032            uc=2.296962e-010 wuc=-3.5392448e-017            vsat=149989.66                  a0=16.704177 la0=-8.5589144e-007            wa0=-1.4731751e-005            pa0=4.9811445e-013 ags=3                          lags=0                          wags=0 pags=0                          keta=0.032837105                lketa=-5.7610972e-009 wketa=-3.6337604e-007            pketa=1.4040829e-014             pclm=1.7105473 lpclm=-3.323244e-008             wpclm=-8.9542246e-007            ppclm=3.6712321e-014 pdiblc2=0.0025559259               lpdiblc2=0                          wpdiblc2=-5.0366889e-010 ppdiblc2=0                          aigbacc=0.0114824                  laigbacc=4.5190832e-011 waigbacc=-1.1286114e-009            paigbacc=5.2446733e-017             aigc=0.010674868 laigc=-2.8334107e-012            waigc=-1.2858253e-011            paigc=2.5478035e-020 aigsd=0.0096513698               laigsd=3.1465495e-012             waigsd=3.2033673e-011 paigsd=-8.0776237e-019            tvoff=0.00231897                 ltvoff=-4.35294e-011 wtvoff=-2.8924e-010               ptvoff=6.75438e-018               kt1=-0.18322836 lkt1=1.329517e-009              wkt1=4.0252512e-008             pkt1=-1.2393462e-015 kt2=-0.058328477               lkt2=-5.3488733e-011            wkt2=-1.5052054e-008 pkt2=4.816657e-016              ute=-0.70403677                lute=-8.1552662e-009 wute=-1.7312354e-007            pute=4.4935984e-015             ua1=1.1116758e-009 lua1=-1.7388961e-017            wua1=-2.8012469e-016            pua1=6.0040425e-024 ub1=8.605396e-019              lub1=-5.0125596e-026            wub1=-2.1542976e-024 pub1=7.1256512e-032             uc1=2.6342848e-010             luc1=-4.0204431e-018 wuc1=-1.6296487e-016            puc1=4.6991188e-024             at=71222.503 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=8.3424289e-010             petab=6.2797849e-018             lu0=-4.627789e-011 pu0=-1.2965897e-017            luc=5.6050078e-019             puc=-3.2513757e-024 lat=0.00028546469              wat=-0.0058158859              pat=1.5728523e-010 lvsat=-0.00038587249             wvsat=-0.045415557               pvsat=1.6359038e-009 leta0=1.3063551e-009             peta0=-6.0559894e-016            eta0_mc=-0.000397205 weta0_mc=3.5812e-09                 u0_sf=-3.97646e-05               wu0_sf=3.5816e-10 vsat_fs=-4667.39                   vsat_ff=-9111.13                   vsat_ss=20260.2 vsat_mc=-397.205                   lu0_sf=1.63035e-12                pu0_sf=-1.46846e-17 lvsat_fs=0.000145778                lvsat_ff=0.000291556                lvsat_ss=-0.000648326 lvsat_mc=1.62854e-05                wvsat_fs=0.00100733                 wvsat_ff=-2.4e-09 wvsat_ss=-0.0183557                 wvsat_mc=0.0035812                  pvsat_fs=3.6e-16 pvsat_ff=2.8e-16                    pvsat_ss=5.87382e-10                pvsat_mc=-1.46829e-10 leta0_mc=1.62854e-11                peta0_mc=-1.46829e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_lvt_mac.8 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=0.3633846 lvth0=2.2140636e-008             wvth0=-2.2090715e-008            pvth0=-3.1919959e-015 k2=-0.0011891992              lk2=-5.2867041e-016            wk2=9.0119658e-010 pk2=2.6800744e-022             cit=0.0040789983               lcit=-5.9072191e-010 wcit=-1.1007708e-009            pcit=1.3411598e-017             voff=-0.15584827 lvoff=-2.1474976e-008            wvoff=3.0727661e-009             pvoff=4.2272704e-016 eta0=-0.0025833333              weta0=6.8705e-009                etab=-0.025989867 wetab=-8.9976068e-009            u0=0.018267222                wu0=7.8082408e-010 ua=-1.3871842e-009            lua=-7.7349308e-017            wua=-4.7730418e-017 pua=3.0019021e-023             ub=1.8408685e-018             wub=3.0199695e-026 uc=1.0750848e-010             wuc=-5.5990044e-018            vsat=120000 a0=2.2238052                  la0=-6.3698905e-007            wa0=5.5477116e-007 pa0=3.4779803e-013             ags=1.3450472                  lags=2.4467451e-007 wags=-7.755862e-008             pags=2.1920457e-013             keta=-0.040621842 lketa=-2.2201861e-008            wketa=8.5585934e-009             pketa=-1.2698356e-014 pclm=0.37520329                 lpclm=2.2307118e-007             wpclm=-7.5999605e-009 ppclm=6.8369245e-014             pdiblc2=0.0014206573               lpdiblc2=7.137668e-010 wpdiblc2=-3.6001438e-012            ppdiblc2=3.2386894e-017             aigbacc=0.013310817 laigbacc=6.4230113e-011             waigbacc=4.0345944e-011             paigbacc=-5.135214e-018 aigc=0.010868708                laigc=-9.9425223e-011            waigc=-3.9113674e-011 paigc=4.874522e-017              aigsd=0.0097002184               laigsd=2.1819645e-010 waigsd=2.8373871e-011             paigsd=-1.3342266e-016            tvoff=0.00166567 ltvoff=-3.70634e-010              wtvoff=4.59336e-011               ptvoff=2.02353e-016 kt1=-0.17707631                lkt1=8.7613073e-012             wkt1=1.280729e-008 pkt1=-6.0985366e-018            kt2=-0.077064895               lkt2=-6.4393768e-013 wkt2=8.0768951e-009             pkt2=5.8250596e-019             ute=-0.9487785 wute=-9.604959e-009             ua1=1.6193134e-009             lua1=-1.61749e-016 wua1=-1.2491512e-016            pua1=1.3482415e-022             ub1=-9.0266023e-019 lub1=-2.5779195e-026            wub1=2.6656541e-026             pub1=-9.058996e-032 uc1=2.6718084e-010             luc1=-1.2817057e-016            wuc1=-8.4245562e-017 puc1=6.5634475e-023             at=140000                     jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)' jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                lu0=0 pu0=0                          luc=1.0564784e-023             puc=-9.5716943e-030 lat=0                          wat=0                          pat=0 lvsat=0                          wvsat=0                          pvsat=0 leta0=0                          peta0=0                          ags_ff=0.222121 ags_fs=0.166591                   ags_ss=0.0573811                  ags_sf=-0.0268397 lags_ff=-1.9902e-07                lags_fs=-1.49266e-07               lags_ss=-5.14133e-08 lags_sf=2.40486e-08                wags_ff=9e-14                      wags_fs=7e-14 wags_ss=-1.52608e-07               wags_sf=-7.63041e-08               pags_ff=3.8e-19 pags_fs=-2.1e-19                   pags_ss=1.36737e-13                pags_sf=6.83682e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.9 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.37914955 lvth0=8.0152459e-009             wvth0=-3.0643355e-008            pvth0=4.4711692e-015 k2=0.0025449072               lk2=-3.3457598e-009            wk2=2.389705e-009 pk2=-1.3337033e-015            cit=0.0057004867               lcit=-2.0435756e-009 wcit=-2.8742246e-009            pcit=1.6024262e-015             voff=-0.17866553 lvoff=-1.0307106e-009            wvoff=5.5986892e-009             pvoff=-1.8405001e-015 eta0=-0.0025833333              weta0=6.8705e-009                etab=-0.025989327 wetab=-8.9979064e-009            u0=0.018213409                wu0=8.1472414e-010 ua=-1.486842e-009             lua=1.1944016e-017             wua=3.003612e-017 pua=-3.9659798e-023            ub=1.8999938e-018             lub=-5.2976309e-026 wub=2.5998277e-026             pub=3.7644702e-033             uc=1.1303811e-010 wuc=-9.4501417e-019            vsat=120000                     a0=1.4206154 la0=8.2668989e-008             wa0=1.4494192e-006             pa0=-4.5380661e-013 ags=1.319744                   lags=2.6734616e-007             wags=-1.1553669e-007 pags=2.5323292e-013             keta=-0.058244132               lketa=-6.4122897e-009 wketa=-1.6310899e-009            pketa=-3.5683995e-015            pclm=0.54900741 lpclm=6.7342696e-008             wpclm=1.3679929e-007             ppclm=-6.1012483e-014 pdiblc2=0.0020361683               lpdiblc2=1.6226892e-010             wpdiblc2=6.4802589e-011 ppdiblc2=-2.8901955e-017            aigbacc=0.01339005                 laigbacc=-6.7633069e-012 waigbacc=-1.3858301e-010            paigbacc=1.5518513e-016             aigc=0.010763483 laigc=-5.1437743e-012            waigc=6.7152263e-011             paigc=-4.6469059e-017 aigsd=0.010148834                laigsd=-1.8376299e-010            waigsd=-2.5949218e-010 paigsd=1.2450532e-016             tvoff=0.00105033                 ltvoff=1.80716e-010 wtvoff=4.27741e-010               ptvoff=-1.39746e-016              kt1=-0.20470127 lkt1=2.476073e-008              wkt1=2.8263743e-008             pkt1=-1.3855081e-014 kt2=-0.08995669                lkt2=1.1550405e-008             wkt2=1.678761e-008 pkt2=-7.8042177e-015            ute=-0.98641347                lute=3.3720929e-008 wute=6.6392217e-008             pute=-6.809347e-014             ua1=1.7179926e-009 lua1=-2.5016554e-016            wua1=1.6842191e-017             pua1=7.8095978e-024 ub1=-7.9380261e-019            lub1=-1.2331563e-025            wub1=-9.0116141e-026 pub1=1.4038362e-032             uc1=1.3842588e-010             luc1=-1.2806125e-017 wuc1=-2.3911308e-018            puc1=-7.7070956e-024            at=98015.311 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-4.8368337e-013            petab=2.6845492e-019             lu0=4.821666e-011 pu0=-3.0374454e-017            luc=-4.9545423e-018            puc=-4.1699848e-024 lat=0.037618281                wat=0.033548395                pat=-3.0059362e-008 lvsat=0                          wvsat=0                          pvsat=0 leta0=0                          peta0=0                          a0_ff=-0.19492 a0_ss=0.495557                   a0_fs=-0.147015                  a0_sf=0.946513 la0_ff=1.74642e-07                la0_ss=-4.44013e-07               la0_fs=1.31725e-07 la0_sf=-8.48069e-07               wa0_ff=-2.72377e-07               wa0_ss=-1.1e-13 wa0_fs=-1.36188e-07               wa0_sf=-4.08566e-07               pa0_ff=2.4405e-13 pa0_ss=1.7e-19                    pa0_fs=1.22025e-13                pa0_sf=3.66075e-13 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.10 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.40917191 lvth0=-5.3747302e-009            wvth0=-2.5983126e-008            pvth0=2.3927075e-015 k2=0.0018601999               lk2=-3.0403804e-009            wk2=5.4569227e-010 pk2=-5.1127358e-016            cit=-8.9099272e-005            lcit=5.385798e-010 wcit=1.3354595e-009             pcit=-2.7509293e-016            voff=-0.18010376 lvoff=-3.8925975e-010            wvoff=4.1798621e-009             pvoff=-1.2077032e-015 eta0=-0.0025833333              weta0=6.8705e-009                etab=-0.016690537 wetab=-1.4075037e-008            u0=0.018069515                wu0=8.0657241e-010 ua=-1.357692e-009             lua=-4.5656867e-017            wua=-6.4383401e-017 pua=2.4513087e-024             ub=1.8158307e-018             lub=-1.5439556e-026 wub=2.099704e-026              pub=5.995022e-033              uc=1.2429659e-010 wuc=-1.560717e-017             vsat=120000                     a0=1.5715803 la0=1.5338678e-008             wa0=8.7980492e-007             pa0=-1.9975865e-013 ags=2.7817718                  lags=-3.847182e-007             wags=-2.765259e-007 pags=3.2503411e-013             keta=-0.04239788                lketa=-1.3479718e-008 wketa=-3.551416e-008             pketa=1.154345e-014              pclm=0.58548374 lpclm=5.1074251e-008             wpclm=1.959759e-009              ppclm=-8.7405251e-016 pdiblc2=0.0018817244               lpdiblc2=2.3115094e-010             wpdiblc2=3.3042866e-010 ppdiblc2=-1.4737118e-016            aigbacc=0.012772954                laigbacc=2.6846145e-010 waigbacc=6.3031061e-010             paigbacc=-1.8774143e-016            aigc=0.010749423 laigc=1.1270693e-012             waigc=-3.6522811e-011            paigc=-2.2997641e-019 aigsd=0.0095602136               laigsd=7.8761639e-011             waigsd=1.4766692e-010 paigsd=-5.7087641e-017            tvoff=0.00175193                 ltvoff=-1.32199e-010 wtvoff=1.12491e-011               ptvoff=4.60093e-017               kt1=-0.13923954 lkt1=-4.435202e-009             wkt1=-5.7171664e-009            pkt1=1.300405e-015 kt2=-0.053034706               lkt2=-4.9168005e-009            wkt2=-4.4348303e-009 pkt2=1.6609905e-015             ute=-0.63176266                lute=-1.2445333e-007 wute=-1.9483113e-007            pute=4.8412145e-014             ua1=1.6577144e-009 lua1=-2.2328145e-016            wua1=2.8127944e-017             pua1=2.7761518e-024 ub1=-1.412911e-018             lub1=1.5280669e-025             wub1=-1.1449724e-025 pub1=2.4912331e-032             uc1=1.0389552e-010             luc1=2.5944159e-018 wuc1=-2.7534472e-017            puc1=3.5068344e-024             at=278306.09 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-4.1477438e-009            petab=2.2646686e-015             lu0=1.1239349e-010 pu0=-2.6738783e-017            luc=-9.9758234e-018            puc=2.3693367e-024 lat=-0.042791407               wat=-0.064959524               pat=1.387517e-008 lvsat=0                          wvsat=0                          pvsat=0 leta0=0                          peta0=0                          vsat_ff=890.881 vsat_ss=-2717.95                   vsat_fs=1811.96                    vsat_sf=-1811.96 a0_ff=0.10607                    a0_ss=-0.568701                  a0_fs=0.0109292 a0_sf=-1.77642                   la0_ff=4.04064e-08                la0_ss=3.06424e-08 la0_fs=6.12829e-08                la0_sf=3.66356e-07                wa0_ff=2.74811e-07 wa0_ss=6.22491e-08                wa0_fs=2.61901e-07                wa0_sf=9.10201e-07 pa0_ff=2.8e-19                    pa0_ss=-2.77617e-14               pa0_fs=-5.55229e-14 pa0_sf=-2.22092e-13               lvsat_ff=-0.00039733                lvsat_ss=0.00121221 lvsat_fs=-0.000808136               lvsat_sf=0.000808136                wvsat_ff=0.00124491 wvsat_ss=-3.3e-09                   wvsat_fs=2.2e-09                    wvsat_sf=-2.2e-09 pvsat_ff=-5.55226e-10               pvsat_ss=1.1e-15                    pvsat_fs=-7e-16 pvsat_sf=7e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.11 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=0.39288203 lvth0=-1.9212746e-009            wvth0=-1.5279549e-008            pvth0=1.2354904e-016 k2=-0.0096454632              lk2=-6.0117983e-010            wk2=-4.2056333e-009 pk2=4.9600742e-016             cit=0.0017033553               lcit=1.5857943e-010 wcit=1.6374819e-010             pcit=-2.669014e-017             voff=-0.17402815 lvoff=-1.6772903e-009            wvoff=-5.9899423e-010            pvoff=-1.9458566e-016 eta0=-0.0025833333              weta0=6.8705e-009                etab=-0.034883666 wetab=2.501849e-009              u0=0.018490559                wu0=8.6920523e-010 ua=-1.7104211e-009            lua=2.9121709e-017             wua=-1.9699412e-018 pua=-1.0780345e-023            ub=1.8294891e-018             lub=-1.8335132e-026 wub=4.5520999e-026             pub=7.9594269e-034             uc=6.51829e-011 wuc=6.0213656e-018             vsat=130717.08                  a0=4.1600718 la0=-5.3342153e-007            wa0=1.7551058e-007             pa0=-5.0448246e-014 ags=-0.10994098                lags=2.283249e-007              wags=1.8330066e-006 pags=-1.2218677e-013            keta=-0.0380561                 lketa=-1.4400175e-008 wketa=3.7243638e-009             pketa=3.2248827e-015             pclm=0.35514165 lpclm=9.9906775e-008             wpclm=1.1443926e-007             ppclm=-2.4719707e-014 pdiblc2=0.0034990199               lpdiblc2=-1.1171571e-010            wpdiblc2=-6.1365323e-010 ppdiblc2=5.2774178e-017             aigbacc=0.015680278                laigbacc=-3.4789112e-010 waigbacc=-1.5154555e-009            paigbacc=2.6716099e-016             aigc=0.010812502 laigc=-1.2245554e-011            waigc=-6.9109982e-011            paigc=6.6785039e-018 aigsd=0.010008067                laigsd=-1.618318e-011             waigsd=-1.1296569e-010 paigsd=-1.8335276e-018            tvoff=0.000613685                ltvoff=1.09109e-010 wtvoff=5.05247e-010               ptvoff=-5.87182e-017              kt1=-0.18748779 lkt1=5.7934261e-009             wkt1=8.0835858e-009             pkt1=-1.6253545e-015 kt2=-0.081716626               lkt2=1.1637665e-009             wkt2=6.0059782e-009 pkt2=-5.5246093e-016            ute=-1.2205936                 lute=3.7882647e-010 wute=2.873314e-008              pute=1.0165188e-015             ua1=1.3901404e-009 lua1=-1.6655576e-016            wua1=-3.675605e-016             pua1=8.6662102e-023 ub1=-1.6281285e-018            lub1=1.9843281e-025             wub1=6.0736219e-025 pub1=-1.2812187e-031            uc1=5.8344974e-011             luc1=1.2251132e-017 wuc1=2.6522311e-017             puc1=-7.9532036e-024            at=100543.36 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-2.9080059e-010            petab=-1.2496312e-015            lu0=2.313212e-011 pu0=-4.0016941e-017            luc=2.5562788e-018             puc=-2.2159128e-024 lat=-0.0051057073              wat=-0.0064891398              pat=1.4794486e-009 lvsat=-0.0022720212              wvsat=-0.0047806613              pvsat=1.0135002e-009 leta0=0                          peta0=0                          vsat_ff=-1654.52 vsat_ss=3329.92                    vsat_fs=-3365.08                   vsat_sf=3365.08 a0_ff=0.689693                   a0_ss=-0.713682                  a0_fs=0.81532 a0_sf=-0.0813224                 la0_ff=-8.33223e-08               la0_ss=6.13764e-08 la0_fs=-1.09247e-07               la0_sf=6.99372e-09                wa0_ff=2.27925e-07 wa0_ss=-1.15598e-07               wa0_fs=-2.81363e-07               wa0_sf=-2.31197e-07 pa0_ff=9.94143e-15                pa0_ss=9.94155e-15                pa0_fs=5.9649e-14 pa0_sf=1.9883e-14                 lvsat_ff=0.000142287                lvsat_ss=-6.99343e-05 lvsat_fs=0.000289396                lvsat_sf=-0.000289396               wvsat_ff=-0.00231198 wvsat_ss=0.000937881                wvsat_fs=4.4e-09                    wvsat_sf=-4.4e-09 pvsat_ff=1.9883e-10                 pvsat_ss=-1.9883e-10                pvsat_fs=1.8e-16 pvsat_sf=-1.8e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.12 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.36178999 lvth0=7.5264023e-010             wvth0=-1.0755898e-008            pvth0=-2.6548492e-016 k2=-0.029686718               lk2=1.1223681e-009             wk2=1.0795168e-008 pk2=-7.9406148e-016            cit=0.0015901957               lcit=1.6831116e-010 wcit=-1.6837617e-010            pcit=1.8725548e-018             voff=-0.17428376 lvoff=-1.6553073e-009            wvoff=-6.4160924e-009            pvoff=3.0568478e-016 eta0=-0.04270272                weta0=2.7821332e-008             etab=-0.077773303 wetab=-1.15073e-008              u0=0.019569245                wu0=4.1274345e-010 ua=-1.4045477e-009            lua=2.8165888e-018             wua=-2.6363885e-016 pua=1.1723181e-023             ub=1.5389487e-018             lub=6.65134e-027 wub=1.7372137e-025             pub=-1.0229289e-032            uc=6.8581362e-011 wuc=-1.462627e-017             vsat=56526.447                  a0=-5.1571575 la0=2.678602e-007              wa0=4.0548308e-006             pa0=-3.8406978e-013 ags=1.913055                   lags=5.4347252e-008             wags=9.8477199e-007 pags=-4.92386e-014              keta=-0.21259574                lketa=6.102337e-010 wketa=1.4763941e-008             pketa=2.2754791e-015             pclm=2.6559897 lpclm=-9.7966156e-008            wpclm=-7.9497036e-007            ppclm=5.3489521e-014 pdiblc2=0.0024777778               lpdiblc2=-2.3888889e-011            wpdiblc2=0 ppdiblc2=0                          aigbacc=0.0083340927               laigbacc=2.8388081e-010 waigbacc=4.9123318e-009             paigbacc=-2.8562872e-016            aigc=0.010715811 laigc=-3.930156e-012             waigc=2.298864e-011              paigc=-1.2419776e-018 aigsd=0.0098685366               laigsd=-4.1836046e-012            waigsd=-1.8319996e-010 paigsd=4.2066196e-018             tvoff=0.00194962                 ltvoff=-5.78168e-012 wtvoff=1.82548e-012               ptvoff=-1.5424e-017               kt1=-0.16886917 lkt1=4.1922255e-009             wkt1=1.1416653e-008             pkt1=-1.9119982e-015 kt2=-0.084196161               lkt2=1.3770066e-009             wkt2=1.5373219e-009 pkt2=-1.6815649e-016            ute=-1.6230976                 lute=3.4994167e-008 wute=1.5083671e-007             pute=-9.4843884e-015            ua1=-9.6630608e-010 lua1=3.6098638e-017             wua1=1.0330167e-015             pua1=-3.3787532e-023 ub1=1.2065383e-018             lub1=-4.5348532e-026            wub1=-1.4218547e-024 pub1=4.6390786e-032             uc1=2.4024444e-010             luc1=-3.3922222e-018 wuc1=-1.1176013e-016            puc1=3.9390867e-024             at=7458.9298 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=3.3977082e-009             petab=-4.4844368e-017            lu0=-6.9634881e-011 pu0=-7.612285e-019             luc=2.264011e-018              puc=-4.4021616e-025 lat=0.0028995535               wat=0.019868543                pat=-7.8731215e-010 lvsat=0.0041083733               wvsat=0.02437116                 pvsat=-1.4935564e-009 leta0=3.4502672e-009             peta0=-1.8017715e-015            vsat_ff=6990.74 vsat_ss=6012.04                    a0_ff=-0.666898                  a0_fs=-1.08694 la0_ff=3.33449e-08                la0_fs=5.43472e-08                wa0_ff=8.20643e-07 wa0_fs=9.84772e-07                pa0_ff=-4.10321e-14               pa0_fs=-4.92386e-14 lvsat_ff=-0.000601204               lvsat_ss=-0.000300602               wvsat_ff=-0.00381694 wvsat_ss=-0.00328257                pvsat_ff=3.28257e-10                pvsat_ss=1.64129e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.13 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.33236571 lvth0=2.2238544e-009             wvth0=2.4711488e-008             pvth0=-2.0388542e-015 k2=-0.059695506               lk2=2.6228075e-009             wk2=2.2818796e-008 pk2=-1.3952429e-015            cit=0.0018394582               lcit=1.5584803e-010 wcit=-8.7302142e-010            pcit=3.7104817e-017             voff=-0.19533283 lvoff=-6.0285374e-010            wvoff=1.4432658e-008             pvoff=-7.3675274e-016 eta0=0.029493449                weta0=-2.3023524e-008            etab=0.031306775 wetab=-5.7409916e-008            u0=0.020218158                wu0=-2.3584655e-010 ua=-1.593854e-009             lua=1.2281908e-017             wua=-2.2879225e-016 pua=9.9808515e-024             ub=1.7479727e-018             lub=-3.799858e-027 wub=8.4986061e-026             pub=-5.7925238e-033            uc=-4.8610253e-011 wuc=5.0139112e-018             vsat=180022.96                  a0=35.348415 la0=-1.7574184e-006            wa0=-2.2185059e-005            pa0=9.279247e-013 ags=3.1229848                  lags=-6.1492407e-009            wags=-1.1142424e-007 pags=5.5712121e-015             keta=-0.44320477                lketa=1.2140685e-008 wketa=2.674698e-007              pketa=-1.0359814e-014            pclm=1.8431471 lpclm=-5.7324028e-008            wpclm=-3.5115833e-007            ppclm=3.1298919e-014 pdiblc2=0.002                      lpdiblc2=0                          wpdiblc2=0 ppdiblc2=0                          aigbacc=0.020784031                laigbacc=-3.3861608e-010 waigbacc=-5.3773896e-009            paigbacc=2.2885735e-016             aigc=0.011038412 laigc=-2.0060207e-011            waigc=-1.8823675e-010            paigc=9.319292e-018 aigsd=0.0096637165               laigsd=6.0573989e-012             waigsd=-2.6257069e-010 paigsd=8.175156e-018              tvoff=0.00785362                 ltvoff=-3.00982e-010 wtvoff=-4.20999e-009              ptvoff=1.95167e-016               kt1=0.32611303 lkt1=-2.0556885e-008            wkt1=-2.9569524e-007            pkt1=1.3443596e-014 kt2=0.012574429                lkt2=-3.4615229e-009            wkt2=-4.5526834e-008 pkt2=2.1850513e-015             ute=-1.1185127                 lute=9.7649266e-009 wute=1.6683159e-007             pute=-1.0284132e-014            ua1=-5.2879592e-009 lua1=2.521813e-016              wua1=3.3171311e-015             pua1=-1.4799325e-022 ub1=6.7298967e-018             lub1=-3.2151646e-025            wub1=-3.9432488e-024 pub1=1.7246049e-031             uc1=3.9228148e-010             luc1=-1.0994074e-017 wuc1=-1.3313502e-016            puc1=5.0078311e-024             at=-53663.156 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-2.0562957e-009            petab=2.2502864e-015             lu0=-1.0208051e-010 pu0=3.1668272e-017             luc=8.1235917e-018             puc=-1.4222252e-024 lat=0.0059556578               wat=0.087274819                pat=-4.157626e-009 lvsat=-0.0020664524              wvsat=-0.050650317               pvsat=2.2575174e-009 leta0=-1.595412e-010             peta0=7.4047127e-016             vsat_ff=-5033.37 lvsat_ff=-1.5e-09                   wvsat_ff=0.00274822                 pvsat_ff=-1.1e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.14 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=0.4220052 lvth0=-1.4513647e-009            wvth0=-4.2081818e-008            pvth0=6.9967133e-016 k2=0.024801265                lk2=-8.4156012e-010            wk2=-6.5832838e-009 pk2=-1.8975761e-016            cit=-0.0077949624              lcit=5.5085927e-010 wcit=3.0180908e-009             pcit=-1.2243078e-016            voff=-0.12364579 lvoff=-3.5420223e-009            wvoff=-1.3537931e-008            pvoff=4.1004141e-016 eta0=0.027903356                weta0=-2.1144651e-008            etab=-0.038099668 wetab=-3.6696617e-009            u0=0.01961227                 wu0=1.6862375e-010 ua=-1.9026312e-009            lua=2.4941773e-017             wua=2.5879016e-016 pua=-1.0010027e-023            ub=1.9719289e-018             lub=-1.2982061e-026 wub=-1.8704459e-025            pub=5.360733e-033              uc=1.2413756e-010 wuc=6.0243682e-017             vsat=108426.78                  a0=-5.0209295 la0=-1.0227531e-007            wa0=4.9511962e-006             pa0=-1.8466176e-013 ags=2.8770152                  lags=3.9355141e-009             wags=1.1142424e-007 pags=-3.5655757e-015            keta=-0.33320974                lketa=7.630889e-009 wketa=-3.1737593e-008            pketa=1.9076892e-015             pclm=-1.6741107 lpclm=8.6883544e-008             wpclm=2.1710777e-006             ppclm=-7.211276e-014 pdiblc2=0.002                      lpdiblc2=0                          wpdiblc2=0 ppdiblc2=0                          aigbacc=0.0035157554               laigbacc=3.693832e-010 waigbacc=6.089169e-009              paigbacc=-2.4127155e-016            aigc=0.01054301 laigc=2.5127861e-013             waigc=1.0660575e-010             paigc=-2.7692505e-018 aigsd=0.0097158109               laigsd=3.9215283e-012             waigsd=-2.6349977e-011 paigsd=-1.5098931e-018            tvoff=0.000468271                ltvoff=1.8177e-012 wtvoff=1.3875e-009                ptvoff=-3.43301e-017              kt1=-0.22394615 lkt1=1.9955414e-009             wkt1=7.7142826e-008             pkt1=-1.8427643e-015 kt2=-0.089406589               lkt2=7.1969881e-010             wkt2=1.3104715e-008 pkt2=-2.1884222e-016            ute=-0.76189928                lute=-4.8562248e-009 wute=-1.207001e-007             pute=1.504667e-015              ua1=1.9898632e-009 lua1=-4.6209425e-017            wua1=-1.0757625e-015            pua1=3.2115383e-023 ub1=-3.98996e-018              lub1=1.1799767e-025             wub1=2.2402551e-024 pub1=-8.1063168e-032            uc1=-3.3733333e-011            luc1=6.4725333e-018 wuc1=1.0626373e-016             puc1=-4.8075179e-024            at=140443.81 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=7.8936849e-010             petab=4.6935997e-017             lu0=-7.7239134e-011 pu0=1.508499e-017              luc=1.0409314e-018             puc=-3.6866458e-024 lat=-0.0020027277              wat=-0.068530389               pat=2.2303876e-009 lvsat=0.00086899116              wvsat=-0.0077595827              pvsat=4.9899732e-010 leta0=-9.4347378e-011            peta0=6.6343747e-016             voff_mc=0.0161778 lvoff_mc=-6.63289e-10               wvoff_mc=-1.46571e-08               pvoff_mc=6.0094e-16 eta0_mc=0.00894815                 weta0_mc=-4.88569e-09               u0_sf=0.000355556 u0_fs=0.000539259                wu0_sf=-1.1e-16                   wu0_fs=-4.88569e-10 vsat_fs=-6251.85                   vsat_ff=-22929.6                   vsat_mc=859.261 lu0_sf=-1.45778e-11               lu0_fs=-2.21096e-11               pu0_sf=-2.4e-23 pu0_fs=2.00313e-17                lvsat_fs=0.000256326                lvsat_ff=0.000733748 lvsat_mc=-3.52296e-05               wvsat_fs=0.00244285                 wvsat_ff=0.0125196 wvsat_mc=0.00244284                 pvsat_fs=-1.00156e-10               pvsat_ff=-4.00626e-10 pvsat_mc=-1.00157e-10               leta0_mc=-3.66874e-10               peta0_mc=2.00313e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.15 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.34309657 lvth0=2.1385251e-008             wvth0=-1.101345e-008             pvth0=-2.779556e-015 k2=-0.00059733221             lk2=5.0652627e-014             wk2=5.7803721e-010 pk2=-2.7676981e-020            cit=0.0016600716               lcit=-6.203682e-010 wcit=2.1996315e-010             pcit=2.9598474e-017             voff=-0.15406802 lvoff=-2.8377233e-008            wvoff=2.100749e-009              pvoff=4.1913592e-015 eta0=0.01277288                 weta0=-1.5139925e-009            etab=-0.043967578 wetab=8.1822347e-010             u0=0.019375803                wu0=1.7553907e-010 ua=-1.5073688e-009            lua=3.4957474e-017             wua=1.7890341e-017 pua=-3.1300482e-023            ub=1.8961623e-018             lub=-7.7188587e-027 wub=9.2764902e-030             pub=4.2144968e-033             uc=1.194898e-010 wuc=-1.2140805e-017            vsat=109777.78                  a0=3.6444039 la0=2.8276691e-012             wa0=-2.2087574e-007            pa0=4.609868e-019 ags=1.261273                   lags=7.4355008e-007             wags=-3.1817902e-008 pags=-5.3181492e-014            keta=-0.033285257               lketa=-5.1829639e-008 wketa=4.552818e-009              pketa=3.478411e-015              pclm=0.35563018 lpclm=3.9915092e-007             wpclm=3.0869597e-009             ppclm=-2.7770289e-014 pdiblc2=0.0014129753               lpdiblc2=7.8287446e-010             wpdiblc2=5.9425208e-013 ppdiblc2=-5.3458918e-018            aigbacc=0.013361814                laigbacc=7.0712616e-011 waigbacc=1.2501119e-011             paigbacc=-8.6746608e-018            aigc=0.010775735 laigc=-9.3383469e-012            waigc=1.1649902e-011             paigc=-4.4221409e-019 aigsd=0.0097760681               laigsd=-1.0952934e-010            waigsd=-1.3040059e-011 paigsd=4.5515615e-017             tvoff=0.00166619                 ltvoff=-9.26517e-014 wtvoff=4.56513e-011               ptvoff=3.76565e-020               kt1=-0.14782321 lkt1=-7.0874165e-012            wkt1=-3.1649e-009               pkt1=2.5548666e-018 kt2=-0.060506488               lkt2=7.9849864e-012             wkt2=-9.6399543e-010 pkt2=-4.1288866e-018            ute=-0.96236289                wute=-2.1878827e-009 ua1=1.2176961e-009             lua1=7.6701183e-017             wua1=9.4367954e-017 pua1=4.6303514e-024             ub1=-5.1069956e-019            lub1=-1.3403975e-025 wub1=-1.8735399e-025            pub1=-3.1479695e-032            uc1=1.5295701e-010 luc1=-1.6098718e-017            wuc1=-2.187935e-017             puc1=4.4432463e-024 at=140000                     jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)' jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                lu0=0 pu0=0                          luc=-1.2051925e-023            puc=2.7770289e-030 lat=0                          wat=0                          pat=0 lvsat=0                          wvsat=0.0055813333               pvsat=0 leta0=0                          peta0=0                          ags_ff=0.278884 ags_fs=0.16659                    ags_ss=-0.278884                  ags_sf=-0.16659 lags_ff=-2.49881e-07               lags_fs=-1.49265e-07               lags_ss=2.49881e-07 lags_sf=1.49265e-07                wags_ff=-3.09933e-08               wags_fs=3.6e-14 wags_ss=3.09933e-08                wags_sf=-3.6e-14                   pags_ff=2.77702e-14 pags_fs=-4.3e-20                   pags_ss=-2.77702e-14               pags_sf=4.3e-20 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.16 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.34590712 lvth0=1.8867001e-008             wvth0=-1.2492989e-008            pvth0=-1.4538892e-015 k2=0.0086709609               lk2=-8.30434e-009              wk2=-9.5512035e-010 pk2=1.3736815e-015             cit=-0.00093737977             lcit=1.7069482e-009 wcit=7.5005052e-010             pcit=-4.453598e-016             voff=-0.18697898 lvoff=1.1109894e-009             wvoff=1.0137833e-008             pvoff=-3.0098683e-015 eta0=0.01277288                 weta0=-1.5139925e-009            etab=-0.043967596 wetab=8.1822845e-010             u0=0.01985411                 wu0=-8.1098507e-011 ua=-1.3988372e-009            lua=-6.2286793e-017            wua=-1.8014464e-017 pua=8.7022387e-025             ub=1.9790547e-018             lub=-8.1990465e-026 wub=-1.7168963e-026            pub=1.96062e-032               uc=1.5034607e-010 wuc=-2.1315157e-017            vsat=109777.78                  a0=5.3365377 la0=-1.516149e-006             wa0=-6.8867434e-007            pa0=4.1914801e-013 ags=1.3361517                  lags=6.7645883e-007             wags=-1.2449524e-007 pags=2.9857405e-014             keta=-0.092271014               lketa=1.0215984e-009 wketa=1.6947588e-008             pketa=-7.6273024e-015            pclm=0.98509962 lpclm=-1.648537e-007             wpclm=-1.0130706e-007            ppclm=6.5766752e-014 pdiblc2=0.0022757587               lpdiblc2=9.820505e-012              wpdiblc2=-6.6013752e-011 ppdiblc2=5.433488e-017              aigbacc=0.012923882                laigbacc=4.6310016e-010 waigbacc=1.1594494e-010             paigbacc=-1.0136033e-016            aigc=0.010919954 laigc=-1.3855909e-010            waigc=-1.8280807e-011            paigc=2.6375701e-017 aigsd=0.0095125767               laigsd=1.2655889e-010             waigsd=8.7904183e-011 paigsd=-4.4930426e-017            tvoff=0.00181592                 ltvoff=-1.34251e-010 wtvoff=9.72684e-012               ptvoff=3.2226e-017                kt1=-0.15018228 lkt1=2.1066358e-009             wkt1=-1.5036274e-009            pkt1=-1.4859454e-015 kt2=-0.051239882               lkt2=-8.2948938e-009            wkt2=-4.3517679e-009 pkt2=3.0313153e-015             ute=-0.93298995                lute=-2.6318153e-008 wute=3.7222978e-008             pute=-3.5312131e-014            ua1=1.4549425e-009 lua1=-1.3587161e-016            wua1=1.6046755e-016             pua1=-5.4594884e-023 ub1=-2.4792464e-019            lub1=-3.6948608e-025            wub1=-3.8816551e-025 pub1=1.4844743e-031             uc1=1.7783414e-010             luc1=-3.8388631e-017 wuc1=-2.390804e-017             puc1=6.2609523e-024             at=160053.31 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=1.6162247e-014             petab=-4.4607802e-021            lu0=-4.2856306e-010 pu0=2.2994727e-016             luc=-2.764723e-017             puc=8.2202227e-024 lat=-0.017967766               wat=-0.00032435249             pat=2.9061983e-010 lvsat=0                          wvsat=0.0055813333               pvsat=0 leta0=0                          peta0=0                          a0_ff=-0.693775 a0_ss=0.495552                   a0_fs=-0.599072                  a0_sf=0.400849 la0_ff=6.21621e-07                la0_ss=-4.44018e-07               la0_fs=5.36768e-07 la0_sf=-3.59161e-07               wa0_ff=5e-13                      wa0_ss=7e-14 wa0_fs=1.10635e-07                wa0_sf=-1.10634e-07               pa0_ff=-4.3e-19 pa0_ss=-1.2e-19                   pa0_fs=-9.91286e-14               pa0_sf=9.91284e-14 pdiblc2_ff=5.06568e-05                pdiblc2_fs=-5.06568e-05               lpdiblc2_ff=-4.53885e-11 lpdiblc2_fs=4.53885e-11                wpdiblc2_ff=-2.76586e-11               wpdiblc2_fs=2.76586e-11 ppdiblc2_ff=2.47821e-17                ppdiblc2_fs=-2.47821e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.17 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.39452475 lvth0=-2.8164609e-009            wvth0=-1.7985773e-008            pvth0=9.9589247e-016 k2=0.00035116794              lk2=-4.5937123e-009            wk2=1.3696238e-009 pk2=3.3684563e-016             cit=0.0037674753               lcit=-3.9141716e-010 wcit=-7.7023023e-010            pcit=2.3268541e-016             voff=-0.17437938 lvoff=-4.5084333e-009            wvoff=1.0543493e-009             pvoff=1.0413656e-015 eta0=0.01277288                 weta0=-1.5139925e-009            etab=-0.043967563 wetab=8.1821946e-010             u0=0.01864379                 wu0=4.93018e-010 ua=-1.4034297e-009            lua=-6.0238565e-017            wua=-3.9410634e-017 pua=1.0412916e-023             ub=1.7519967e-018             lub=1.9277403e-026 wub=5.5850402e-026             pub=-1.2960438e-032            uc=1.0956938e-010 wuc=-7.5661143e-018            vsat=109777.78                  a0=2.1593249 la0=-9.9112138e-008            wa0=5.5889631e-007             pa0=-1.372685e-013 ags=1.8611863                  lags=4.4229338e-007             wags=2.2611376e-007 pags=-1.2651421e-013            keta=-0.11033122                lketa=9.0764491e-009 wketa=1.5774419e-009             pketa=-7.7221746e-016            pclm=0.55711194 lpclm=2.6028803e-008             wpclm=1.7450764e-008             ppclm=1.2800762e-014 pdiblc2=0.0023920208               lpdiblc2=-4.2032395e-011            wpdiblc2=5.1806793e-011 ppdiblc2=1.7869171e-018             aigbacc=0.013784604                laigbacc=7.92182e-011 waigbacc=7.7950072e-011             paigbacc=-8.4414614e-017            aigc=0.010595611 laigc=6.0980392e-012             waigc=4.7458716e-011             paigc=-2.944126e-018 aigsd=0.0099325161               laigsd=-6.0734064e-011            waigsd=-5.5610252e-011 paigsd=1.9077012e-017             tvoff=0.00149903                 ltvoff=7.08324e-012 wtvoff=1.49334e-010               ptvoff=-3.00388e-017              kt1=-0.13686655 lkt1=-3.8321778e-009            wkt1=-7.0128184e-009            pkt1=9.7115383e-016 kt2=-0.069691801               lkt2=-6.5337668e-011            wkt2=4.659944e-009 pkt2=-9.8790824e-016            ute=-0.82255519                lute=-7.5572057e-008 wute=-9.0658416e-008            pute=2.1722971e-014             ua1=1.7597317e-009 lua1=-2.718076e-016             wua1=-2.7573509e-017            pua1=2.9271427e-023 ub1=-1.6161115e-018            lub1=2.4072526e-025             wub1=-3.5497271e-027 pub1=-2.3091209e-032            uc1=8.0511573e-011             luc1=5.0172354e-018 wuc1=-1.4766835e-017            puc1=2.1839749e-024             at=155970.58 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=1.6342321e-015             petab=-4.5104806e-022            lu0=1.1123948e-010 pu0=-2.6108691e-017            luc=-9.4608286e-018            puc=2.0881495e-024 lat=-0.016146868               wat=0.0018356653               pat=-6.727481e-010 lvsat=0                          wvsat=0.0055813333               pvsat=0 leta0=0                          peta0=0                          vsat_ff=3170.94 vsat_ss=-2717.95                   vsat_fs=1811.97                    vsat_sf=-1811.97 a0_ff=0.609396                   a0_ss=-0.454701                  a0_fs=0.972878 a0_sf=-0.499069                  la0_ff=4.04069e-08                la0_ss=-2.02038e-08 la0_fs=-1.64321e-07               la0_sf=4.22025e-08                wa0_ff=-4.1e-13 wa0_ss=-4.1e-13                   wa0_fs=-2.63324e-07               wa0_sf=2.12759e-07 pa0_ff=2.2e-19                    pa0_ss=-2.2e-19                   pa0_fs=6.76572e-14 pa0_sf=-4.51048e-14               pdiblc2_ff=-9.74169e-05               pdiblc2_fs=9.74169e-05 lpdiblc2_ff=2.06524e-11                lpdiblc2_fs=-2.06524e-11               wpdiblc2_ff=5.31896e-11 wpdiblc2_fs=-5.31896e-11               ppdiblc2_ff=-1.12762e-17               ppdiblc2_fs=1.12762e-17 lvsat_ff=-0.00141424                lvsat_ss=0.00121221                 lvsat_fs=-0.000808135 lvsat_sf=0.000808135                wvsat_ff=-2.6e-09                   wvsat_ss=2.2e-09 wvsat_fs=-1.5e-09                   wvsat_sf=1.5e-09                    pvsat_ff=-1e-16 pvsat_ss=9e-17                      pvsat_fs=-6e-17                     pvsat_sf=6e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.18 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.39053011 lvth0=-1.9695982e-009            wvth0=-1.3995401e-008            pvth0=1.499337e-016 k2=-0.024015126               lk2=5.7194199e-010             wk2=3.6402026e-009 pk2=-1.4451709e-016            cit=0.00080696852              lcit=2.3621027e-010 wcit=6.5317536e-010             pcit=-6.9076578e-017            voff=-0.19338875 lvoff=-4.7844652e-010            wvoff=9.9718959e-009             pvoff=-8.4915434e-016 eta0=0.014665481                weta0=-2.5473525e-009            etab=-0.029128047 wetab=-6.4071884e-010            u0=0.019620923                wu0=2.5202625e-010 ua=-1.7438712e-009            lua=1.1935036e-017             wua=1.6293787e-017 pua=-1.3964216e-024            ub=1.9623113e-018             lub=-2.5309289e-026 wub=-2.699993e-026             pub=4.6038329e-033             uc=7.1512309e-011 wuc=2.5655083e-018             vsat=107393.11                  a0=4.6200571 la0=-6.2078735e-007            wa0=-7.5641392e-008            pa0=-2.7465066e-015 ags=3.4823844                  lags=9.8599375e-008             wags=-1.2840312e-007 pags=-5.1356634e-014            keta=-0.066750186               lketa=-1.6272944e-010 wketa=1.9391335e-008             pketa=-4.5487628e-015            pclm=0.38109874 lpclm=6.33436e-008               wpclm=1.0026669e-007             ppclm=-4.7562133e-015 pdiblc2=0.0022592629               lpdiblc2=-1.3887723e-011            wpdiblc2=6.3254051e-011 ppdiblc2=-6.3990177e-019            aigbacc=0.012938289                laigbacc=2.5863693e-010 waigbacc=-1.8329596e-011            paigbacc=-6.4003324e-017            aigc=0.010637484 laigc=-2.7790391e-012            waigc=2.6449694e-011             paigc=1.5097866e-018 aigsd=0.0097544161               laigsd=-2.2976864e-011            waigsd=2.552743e-011 paigsd=1.8758238e-018             tvoff=0.0013081                  ltvoff=4.75602e-011 wtvoff=1.26097e-010               ptvoff=-2.51126e-017              kt1=-0.15524715 lkt1=6.4508675e-011             wkt1=-9.5198025e-009            pkt1=1.5026345e-015 kt2=-0.070716665               lkt2=1.5193333e-010             wkt2=-5.5813335e-016 pkt2=5.7930019e-030             ute=-1.189276                  lute=2.172764e-009 wute=1.1633762e-008             pute=3.7028922e-017             ua1=1.7711289e-010 lua1=6.3707594e-017             wua1=2.947525e-016              pua1=-3.9061687e-023 ub1=1.1966885e-019             lub1=-1.2726017e-025            wub1=-3.4693515e-025 pub1=4.97065e-032               uc1=1.5417002e-010             luc1=-1.0598355e-017 wuc1=-2.5798163e-017            puc1=4.5226164e-024             at=91739.933 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-3.1459758e-009            petab=3.0929447e-016             lu0=-9.5912754e-011 pu0=2.498156e-017              luc=-1.3927293e-018            puc=-5.9754431e-026 lat=-0.0025299709              wat=-0.0016824695              pat=7.3096465e-011 lvsat=0.00050554909              wvsat=0.0079542258               pvsat=-5.0305321e-010 leta0=-4.0123135e-010            peta0=2.1907232e-016             vsat_ff=-5888.85 vsat_ss=5047.61                    vsat_fs=-3365.08                   vsat_sf=3365.08 a0_ff=1.10714                    a0_ss=-0.925399                  a0_fs=0.0582357 a0_sf=-0.504761                  la0_ff=-6.51148e-08               la0_ss=7.95843e-08 la0_fs=2.95828e-08                la0_sf=4.34095e-08                wa0_ff=1.5e-13 wa0_ss=1.9e-13                    wa0_fs=1.32003e-07                wa0_sf=-4.4e-13 pa0_ff=-4.7e-20                   pa0_ss=-4.6e-20                   pa0_fs=-1.61522e-14 pa0_sf=2e-21                      lvsat_ff=0.000506441                lvsat_ss=-0.000434095 lvsat_fs=0.000289397                lvsat_sf=-0.000289397               wvsat_ff=4.8e-09 wvsat_ss=4.4e-09                    wvsat_fs=-3e-09                     wvsat_sf=3e-09 pvsat_ff=-4.7e-16                   pvsat_ss=-2e-17                     pvsat_fs=1e-17 pvsat_sf=-1e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.19 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.37218248 lvth0=-3.9170201e-010            wvth0=-1.6430195e-008            pvth0=3.5932594e-016 k2=-0.011028039               lk2=-5.4494747e-010            wk2=6.0752939e-010 pk2=1.1629281e-016             cit=0.0016926013               lcit=1.6004585e-010 wcit=-2.2428962e-010            pcit=6.3854111e-018             voff=-0.18734149 lvoff=-9.9851135e-010            wvoff=7.1342463e-010             pvoff=-5.2925812e-017 eta0=0.010143635                weta0=-1.0327781e-009            etab=-0.11273872 wetab=7.5838189e-009             u0=0.018527944                wu0=9.8129378e-010 ua=-1.8983837e-009            lua=2.522311e-017              wua=5.9956174e-018 pua=-5.1077899e-025            ub=1.8101264e-018             lub=-1.2221384e-026 wub=2.5658385e-026             pub=7.5217831e-035             uc=6.2586295e-011 wuc=-1.1352964e-017            vsat=97514.089                  a0=2.7496256 la0=-4.5993025e-007            wa0=-2.6227283e-007            pa0=1.3303797e-014 ags=5.4714812                  lags=-7.2462951e-008            wags=-9.5812876e-007 pags=1.9999771e-014             keta=-0.067374102               lketa=-1.0907269e-010 wketa=-6.4527074e-008            pketa=2.6682204e-015             pclm=1.0032803 lpclm=9.8359835e-009             wpclm=1.0740894e-007             ppclm=-5.370447e-015 pdiblc2=0.0022335803               lpdiblc2=-1.1679012e-011            wpdiblc2=1.3333185e-010 ppdiblc2=-6.6665926e-018            aigbacc=0.020245742                laigbacc=-3.6980398e-010 waigbacc=-1.5914284e-009            paigbacc=7.1283175e-017             aigc=0.010563019 laigc=3.6249162e-012             waigc=1.0641288e-010             paigc=-5.367047e-018 aigsd=0.0093976694               laigsd=7.703353e-012              waigsd=7.3893512e-011 paigsd=-2.2836593e-018            tvoff=0.00326718                 ltvoff=-1.20921e-010 wtvoff=-7.17561e-010              ptvoff=4.7442e-017                kt1=-0.16221506 lkt1=6.6374919e-010             wkt1=7.783507e-009              pkt1=1.4549838e-017 kt2=-0.095578082               lkt2=2.2900152e-009             wkt2=7.7518505e-009 pkt2=-6.6665919e-016            ute=-1.5197781                 lute=3.0595939e-008 wute=9.4424284e-008             pute=-7.082956e-015             ua1=1.6659065e-009 lua1=-6.432866e-017             wua1=-4.0417144e-016            pua1=2.1045772e-023 ub1=-2.7610445e-018            lub1=1.2048117e-025             wub1=7.4444547e-025 pub1=-4.4152233e-032            uc1=-7.0301235e-011            luc1=8.7061728e-018 wuc1=5.7797807e-017             puc1=-2.666637e-024             at=38972.13 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=4.0445423e-009             petab=-3.9801578e-016            lu0=-1.9165312e-012 pu0=-3.7735447e-017            luc=-6.2509212e-019            puc=1.1372341e-024 lat=0.0020080602               wat=0.0026623359               pat=-3.0055679e-010 lvsat=0.0013551451               wvsat=0.0019919068               pvsat=9.7062255e-012 leta0=-1.2352602e-011            peta0=8.8818913e-017             vsat_ff=-1419.75 a0_ff=0.836109                   a0_fs=0.960865                   la0_ff=-4.18055e-08 la0_fs=-4.80432e-08               wa0_ff=4.8e-13                    wa0_fs=-1.33332e-07 pa0_ff=2.6e-20                    pa0_fs=6.66662e-15                lvsat_ff=0.000122099 wvsat_ff=0.000775185                pvsat_ff=-6.66659e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.20 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.38078395 lvth0=-8.2177556e-010            wvth0=-1.7248705e-009            pvth0=-3.7594027e-016 k2=-0.028714841               lk2=3.3939263e-010             wk2=5.9033534e-009 pk2=-1.4849839e-016            cit=-0.00032615506             lcit=2.6098367e-010 wcit=3.0940344e-010             pcit=-2.0299242e-017            voff=-0.098232489 lvoff=-5.4539611e-009            wvoff=-3.858413e-008             pvoff=1.9119519e-015 eta0=-0.0085471174              weta0=-2.253375e-009             etab=-0.070387499 wetab=-1.8848426e-009            u0=0.019077175                wu0=3.8713015e-010 ua=-1.9395886e-009            lua=2.7283357e-017             wua=-4.0021171e-017 pua=1.7900604e-024             ub=1.8648669e-018             lub=-1.495841e-026 wub=2.1161832e-026             pub=3.0004547e-034             uc=-1.887609e-010 wuc=8.1536166e-017             vsat=34324.986                  a0=-13.623964 la0=3.5874926e-007             wa0=4.5538605e-006             pa0=-2.2750287e-013 ags=3.8582425                  lags=8.1989876e-009             wags=-5.1287492e-007 pags=-2.2629206e-015            keta=0.20681481                 lketa=-1.3818518e-008 wketa=-8.7440889e-008            pketa=3.8139111e-015             pclm=1.2 lpclm=0                          wpclm=0                          ppclm=0 pdiblc2=0.002                      lpdiblc2=0                          wpdiblc2=0 ppdiblc2=0                          aigbacc=0.014013507                laigbacc=-5.8192255e-011 waigbacc=-1.6806837e-009            paigbacc=7.574594e-017              aigc=0.010688217 laigc=-2.6349637e-012            waigc=2.9697531e-012             paigc=-1.9489086e-019 aigsd=0.0089606855               laigsd=2.9552545e-011             waigsd=1.2128421e-010 paigsd=-4.653194e-018             tvoff=-0.00306309                ltvoff=1.95593e-010 wtvoff=1.75054e-009               ptvoff=-7.59628e-017              kt1=-0.44414101 lkt1=1.4760046e-008             wkt1=1.2486346e-007             pkt1=-5.839448e-015 kt2=-0.022747574               lkt2=-1.3515102e-009            wkt2=-2.624102e-008 pkt2=1.0329843e-015             ute=-0.70415475                lute=-1.0185227e-008 wute=-5.9407873e-008            pute=6.086519e-016              ua1=1.4218717e-009 lua1=-5.2126916e-017            wua1=-3.464366e-016             pua1=1.815903e-023 ub1=-9.2541361e-019            lub1=2.869963e-026              wub1=2.3655068e-025 pub1=-1.8757494e-032            uc1=-8.7506173e-012            luc1=5.628642e-018 wuc1=8.5828504e-017             puc1=-4.0681719e-024            at=182610.8 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=1.9269811e-009             petab=7.5417295e-017             lu0=-2.9378059e-011 pu0=-8.0272659e-018            luc=1.1942268e-017             puc=-3.5072223e-024 lat=-0.0051738732              wat=-0.041730759               pat=1.9190979e-009 lvsat=0.0045146002               wvsat=0.028900778                pvsat=-1.3357373e-009 leta0=9.2218501e-010             peta0=1.4984876e-016             vsat_ff=5679.01 vsat_fs=4656.79                    lvsat_ff=-0.00023284                lvsat_fs=-0.00023284 wvsat_ff=-0.00310074                wvsat_fs=-0.00254261                pvsat_ff=1.2713e-10 pvsat_fs=1.2713e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.21 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=0.39141669 lvth0=-1.257718e-009             wvth0=-2.5380493e-008            pvth0=5.9394024e-016 k2=0.005675318                lk2=-1.0706039e-009            wk2=3.8594831e-009 pk2=-6.4699709e-017            cit=0.0067701021               lcit=-2.9962873e-011 wcit=-4.9344344e-009            pcit=1.9469811e-016             voff=-0.20556148 lvoff=-1.0534725e-009            wvoff=3.1188034e-008             pvoff=-9.4870679e-016 eta0=-0.019928499               weta0=4.9715417e-009             etab=-0.039938822 wetab=-2.6654836e-009            u0=0.020028851                wu0=-5.8829548e-011 ua=-1.3447086e-009            lua=2.8932768e-018             wua=-4.5835587e-017 pua=2.0284515e-024             ub=1.4489204e-018             lub=2.0953965e-027 wub=9.8518038e-026             pub=-2.871559e-033             uc=2.178087e-010 wuc=9.0992402e-018             vsat=166649.59                  a0=11.665382 la0=-6.7811396e-007            wa0=-4.1595299e-006            pa0=1.2974614e-013 ags=4.186202                   lags=-5.2473521e-009            wags=-6.0339174e-007 pags=1.4482692e-015             keta=-0.52006558                lketa=1.5983578e-008 wketa=7.0285694e-008             pketa=-2.6528788e-015            pclm=1.7933826 lpclm=-2.4328687e-008            wpclm=2.7782639e-007             ppclm=-1.1390882e-014 pdiblc2=0.002                      lpdiblc2=0                          wpdiblc2=0 ppdiblc2=0                          aigbacc=0.014629558                laigbacc=-8.3450338e-011 waigbacc=2.1032889e-011             paigbacc=5.9755586e-018             aigc=0.01070584 laigc=-3.3575123e-012            waigc=1.7700479e-011             paigc=-7.9885063e-019 aigsd=0.0096267261               laigsd=2.2448825e-012             waigsd=2.2290317e-011 paigsd=-5.9444453e-019            tvoff=0.00309383                 ltvoff=-5.68412e-011 wtvoff=-4.60622e-011              ptvoff=-2.30232e-018              kt1=-0.10131145 lkt1=7.0403452e-010             wkt1=1.0184281e-008             pkt1=-1.1376015e-015 kt2=-0.073249258               lkt2=7.1905886e-010             wkt2=4.2828127e-009 pkt2=-2.184928e-016             ute=-0.93680972                lute=-6.4637348e-010 wute=-2.5199001e-008            pute=-7.9391187e-016            ua1=-4.6009492e-010 lua1=2.5033713e-017             wua1=2.6191464e-016             pua1=-6.7833708e-024 ub1=1.6719823e-018             lub1=-7.7793602e-026            wub1=-8.5116545e-025 pub1=2.5838867e-032             uc1=3.3080494e-010             luc1=-8.2931358e-018 wuc1=-9.2774163e-017            puc1=3.2545375e-024             at=51260.966 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=6.7858537e-010             petab=1.0742358e-016             lu0=-6.8396811e-011 pu0=1.0257082e-017             luc=-4.7270859e-018            puc=-5.3730838e-025 lat=0.00021146988              wat=-0.019836557               pat=1.0214357e-009 lvsat=-0.00091070856             wvsat=-0.039549239               pvsat=1.4707134e-009 leta0=1.3888216e-009             peta0=-1.4637282e-016            cit_mcl=0.00363457 lcit_mcl=-1.49017e-10               wcit_mcl=-1.98447e-09               pcit_mcl=8.13634e-17 voff_ff=0.0181728                  voff_mc=-0.0215704                 lvoff_ff=-7.45086e-10 lvoff_mc=8.84385e-10                wvoff_ff=-9.92237e-09               wvoff_mc=5.95342e-09 pvoff_ff=4.06817e-16                pvoff_mc=-2.4409e-16                u0_sf=0.00144593 u0_fs=-0.000719012               u0_ss=0.00218074                 u0_ff=-0.0012721 wu0_sf=-5.95342e-10               wu0_fs=1.98447e-10                wu0_ss=-1.19068e-09 wu0_ff=6.94566e-10                vsat_fs=-8251.85                   vsat_ss=10903.7 vsat_ff=-14538.3                   vsat_sf=7269.14                    vsat_mc=10785.2 lu0_sf=-5.9283e-11                lu0_fs=2.94795e-11                lu0_ss=-8.94104e-11 lu0_ff=5.2156e-11                 pu0_sf=2.4409e-17                 pu0_fs=-8.13634e-18 pu0_ss=4.88181e-17                pu0_ff=-2.84772e-17               lvsat_fs=0.000296415 lvsat_ss=-0.000447052               lvsat_ff=0.000596069                lvsat_sf=-0.000298035 lvsat_mc=-0.000442193               wvsat_fs=0.00353484                 wvsat_ss=-0.00595342 wvsat_ff=0.0079379                  wvsat_sf=-0.00396895                wvsat_mc=-0.00297671 pvsat_fs=-1.22045e-10               pvsat_ss=2.4409e-10                 pvsat_ff=-3.25454e-10 pvsat_sf=1.62727e-10                pvsat_mc=1.22045e-10 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.22 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.32949898 lvth0=1.6685798e-008             wvth0=-7.2605145e-009            pvth0=-1.4825069e-015 k2=-0.012643196               lk2=-2.3783645e-013            wk2=3.9026956e-009 pk2=5.1946004e-020             cit=0.0026582337               lcit=-4.2391472e-010 wcit=-5.5529596e-011            pcit=-2.4622686e-017            voff=-0.15874432 lvoff=-1.0022904e-008            wvoff=3.3914074e-009             pvoff=-8.7443542e-016 eta0=0.0067859406               weta0=1.3840278e-010             etab=-0.041003 u0=0.019057205                wu0=2.6347216e-010             ua=-1.497928e-009 lua=-2.4829248e-017            wua=1.5284681e-017             pua=-1.4799347e-023 ub=1.7996762e-018             lub=1.2864765e-026             wub=2.6639438e-026 pub=-1.4665831e-033            uc=4.9211413e-011             wuc=7.256029e-018 vsat=125074.07                  a0=2.2347367                  la0=4.0505811e-007 wa0=1.6819242e-007             pa0=-1.117948e-013             ags=0.97536027 lags=5.8704434e-007             wags=4.7094016e-008             pags=-9.9859076e-015 keta=0.014768148                lketa=-4.552642e-008             wketa=-8.7099217e-009 pketa=1.7387224e-015             pclm=0.24861686                 lpclm=9.5739001e-008 wpclm=3.2622635e-008             ppclm=5.5971399e-014             pdiblc2=0.0014565982 lpdiblc2=3.904426e-010              wpdiblc2=-1.1445676e-011            ppdiblc2=1.029653e-016 aigbacc=0.013296543                laigbacc=2.8621295e-011             waigbacc=3.0516055e-011 paigbacc=2.9425439e-018             aigc=0.010758465                laigc=-1.2052102e-011 waigc=1.6416306e-011             paigc=3.0678235e-019             aigsd=0.0096396423 laigsd=1.2822695e-010             waigsd=2.4613446e-011             paigsd=-2.0105122e-017 tvoff=0.0017889                  ltvoff=7.77356e-011               wtvoff=1.17843e-011 ptvoff=-2.14429e-017              kt1=-0.14283744                lkt1=3.276502e-013 wkt1=-4.5409721e-009            pkt1=5.0830819e-019             kt2=-0.062948753 lkt2=-1.1882903e-011            wkt2=-2.8993014e-010            pkt2=1.354651e-018 ute=-0.80864222                wute=-4.4614787e-008            ua1=1.5510458e-009 lua1=1.7051176e-016             wua1=2.3634246e-018             pua1=-2.1261368e-023 ub1=-1.1191418e-018            lub1=-1.4371025e-025            wub1=-1.9423934e-026 pub1=-2.8810638e-032            uc1=6.9267143e-011             luc1=2.9601932e-017 wuc1=1.2190526e-018             puc1=-8.1701332e-024            at=140000 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' lu0=0                          pu0=0                          luc=-3.3907557e-024 puc=3.8654616e-031             lat=0                          wat=0 pat=0                          lvsat=0                          wvsat=0.0013595556 pvsat=0                          leta0=0                          peta0=0 ags_ff=0.127514                   ags_fs=0.166591                   ags_ss=-0.166591 ags_sf=-0.143145                  lags_ff=-1.14253e-07               lags_fs=-1.49266e-07 lags_ss=1.49266e-07                lags_sf=1.28258e-07                wags_ff=1.07852e-08 wags_fs=-1.4e-14                   wags_ss=1.4e-14                    wags_sf=-6.4711e-09 pags_ff=-9.66354e-15               pags_fs=-5e-21                     pags_ss=5e-21 pags_sf=5.79813e-15 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.23 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.32507131 lvth0=2.065299e-008              wvth0=-6.7423056e-009            pvth0=-1.9468221e-015 k2=-0.015378049               lk2=2.4501907e-009             wk2=5.6824064e-009 pk2=-1.594569e-015             cit=0.0020963541               lcit=7.9529421e-011 wcit=-8.7260022e-011            pcit=3.8077752e-018             voff=-0.15715236 lvoff=-1.1449301e-008            wvoff=1.9056849e-009             pvoff=4.5677193e-016 eta0=0.0067859406               weta0=1.3840278e-010             etab=-0.041003 u0=0.018339467                wu0=3.369428e-010              ua=-1.520285e-009 lua=-4.7973437e-018            wua=1.5505125e-017             pua=-1.4996864e-023 ub=1.8074082e-018             lub=5.9369193e-027             wub=3.0205482e-026 pub=-4.6617585e-033            uc=2.8956145e-011             wuc=1.2188461e-017 vsat=125074.07                  a0=2.2023236                  la0=4.3410018e-007 wa0=1.7636872e-007             pa0=-1.1912076e-013            ags=0.51156286 lags=1.0026068e-006             wags=1.0309127e-007             pags=-6.0159443e-014 keta=0.036989699                lketa=-6.543693e-008             wketa=-1.8728369e-008 pketa=1.0715251e-014             pclm=0.13971672                 lpclm=1.9331353e-007 wpclm=1.3201862e-007             ppclm=-3.3087404e-014            pdiblc2=0.0014993559 lpdiblc2=3.5213173e-010             wpdiblc2=1.4827343e-010             ppdiblc2=-4.0143017e-017 aigbacc=0.012887276                laigbacc=3.9532497e-010             waigbacc=1.2604833e-010 paigbacc=-8.2654374e-017            aigc=0.010800202                laigc=-4.944875e-011 waigc=1.4770697e-011             paigc=1.7812484e-018             aigsd=0.0098922388 laigsd=-9.809946e-011             waigsd=-1.6882536e-011            paigsd=1.7075279e-017 tvoff=0.00175793                 ltvoff=1.0548e-010                wtvoff=2.57317e-011 ptvoff=-3.39398e-017              kt1=-0.13642086                lkt1=-5.7489337e-009 wkt1=-5.3017795e-009            pkt1=6.8219182e-016             kt2=-0.068266885 lkt2=4.753163e-009              wkt2=3.476849e-010              pkt2=-5.6994842e-016 ute=-0.5095503                 lute=-2.6798636e-007            wute=-7.9646366e-008 pute=3.1388295e-014             ua1=2.0941047e-009             lua1=-3.1606895e-016 wua1=-1.5941207e-017            pua1=-4.8604184e-024            ub1=-1.3170567e-018 lub1=3.3621487e-026             wub1=-9.308507e-026             pub1=3.7189741e-032 uc1=1.4819843e-010             luc1=-4.1120498e-017            wuc1=-1.5728582e-017 puc1=7.0149477e-024             at=170767.83 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' lu0=6.4309262e-010             pu0=-6.5829696e-017            luc=1.8148717e-017 puc=-4.4194587e-024            lat=-0.027567971               wat=-0.0032815587 pat=2.9402766e-009             lvsat=0                          wvsat=0.0013595556 pvsat=0                          leta0=0                          peta0=0 a0_ff=-0.763521                  a0_ss=0.84428                    a0_fs=-0.337712 la0_ff=6.84112e-07                la0_ss=-7.56475e-07               la0_fs=3.0259e-07 wa0_ff=1.92495e-08                wa0_ss=-9.62479e-08               wa0_fs=3.84992e-08 pa0_ff=-1.72473e-14               pa0_ss=8.62381e-14                pa0_fs=-3.44952e-14 pdiblc2_ff=-4.95556e-05               pdiblc2_fs=4.95556e-05                lpdiblc2_ff=4.44018e-11 lpdiblc2_fs=-4.44018e-11               wpdiblc2_ff=1e-19                      wpdiblc2_fs=-1e-19 ppdiblc2_ff=-2e-24                     ppdiblc2_fs=2e-24 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.24 nmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.37294757 lvth0=-6.9982425e-010            wvth0=-1.2030473e-008            pvth0=4.1170075e-016 k2=0.00036962387              lk2=-4.5732714e-009            wk2=1.3645299e-009 pk2=3.3120395e-016             cit=0.0013100018               lcit=4.3024252e-010 wcit=-9.1967556e-011            pcit=5.9073353e-018             voff=-0.1860512 lvoff=1.4395824e-009             wvoff=4.2757717e-009             pvoff=-6.0028679e-016 eta0=0.0067859406               weta0=1.3840278e-010             etab=-0.041003 u0=0.019699902                wu0=2.0153112e-010             ua=-1.5044092e-009 lua=-1.1877967e-017            wua=-1.154029e-017             pua=-2.934609e-024 ub=1.8754563e-018             lub=-2.4412552e-026            wub=2.1775553e-026 pub=-9.0201004e-034            uc=6.9237193e-011             wuc=3.5655697e-018 vsat=125074.07                  a0=4.6131719                  la0=-6.4113815e-007 wa0=-1.1836545e-007            pa0=1.2330678e-014             ags=3.0246263 lags=-1.1821948e-007            wags=-9.4995686e-008            pags=2.8187337e-014 keta=-0.15285362                lketa=1.9233192e-008             wketa=1.3313626e-008 pketa=-3.5754787e-015            pclm=0.30593866                 lpclm=1.1917854e-007 wpclm=8.677459e-008              ppclm=-1.2908566e-014            pdiblc2=0.0024247194 lpdiblc2=-6.0580394e-011            wpdiblc2=4.2781992e-011             ppdiblc2=6.906165e-018 aigbacc=0.014329725                laigbacc=-2.4800738e-010            waigbacc=-7.2503288e-011 paigbacc=5.8996475e-018             aigc=0.010690869                laigc=-6.8619041e-013 waigc=2.1167394e-011             paigc=-1.0716786e-018            aigsd=0.0096045323 laigsd=3.0217644e-011             waigsd=3.4913288e-011             paigsd=-6.0256589e-018 tvoff=0.00227307                 ltvoff=-1.24271e-010              wtvoff=-6.43016e-011 ptvoff=6.21505e-018               kt1=-0.14156567                lkt1=-3.4543473e-009 wkt1=-5.715862e-009             pkt1=8.6687261e-016             kt2=-0.050049287 lkt2=-3.3718855e-009            wkt2=-7.6138993e-010            pkt2=-7.5301049e-017 ute=-1.1118551                 lute=6.415678e-010              wute=-1.0811646e-008 pute=6.880102e-016              ua1=1.5786903e-009             lua1=-8.6194141e-017 wua1=2.2393923e-017             pua1=-2.1957886e-023            ub1=-1.3149249e-018 lub1=3.2670714e-026             wub1=-8.6677236e-026            pub1=3.4331847e-032 uc1=3.2108895e-011             luc1=1.0655433e-017             wuc1=-1.4076961e-018 puc1=6.2783246e-025             at=151297.53 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' lu0=3.6338737e-011             pu0=-5.4360874e-018            luc=1.8336972e-019 puc=-5.7364919e-025            lat=-0.018884219               wat=0.0031254276 pat=8.2760718e-011             lvsat=0                          wvsat=0.0013595556 pvsat=0                          leta0=0                          peta0=0 vsat_ff=3808.48                    vsat_ss=-4630.58                   vsat_fs=3087.05 vsat_sf=-3087.05                   a0_ff=0.743527                   a0_ss=-0.77468 a0_fs=0.0320354                  a0_sf=0.463058                   la0_ff=1.19725e-08 la0_ss=-3.4421e-08                la0_fs=1.37682e-07                la0_sf=-2.06524e-07 wa0_ff=-3.70176e-08               wa0_ss=8.83129e-08                wa0_fs=-3.652e-09 wa0_sf=-5.27886e-08               pa0_ff=7.84785e-15                pa0_ss=3.92398e-15 pa0_fs=-1.56958e-14               pa0_sf=2.35437e-14                pdiblc2_ff=0.000127176 pdiblc2_fs=-0.000127176               lpdiblc2_ff=-3.44206e-11               lpdiblc2_fs=3.44206e-11 wpdiblc2_ff=-8.7981e-12                wpdiblc2_fs=8.7981e-12                 ppdiblc2_ff=3.92395e-18 ppdiblc2_fs=-3.92395e-18               lvsat_ff=-0.00169858                lvsat_ss=0.00206524 lvsat_fs=-0.00137683                lvsat_sf=0.00137683                 wvsat_ff=-0.000175962 wvsat_ss=0.000527886                wvsat_fs=-0.000351924               wvsat_sf=0.000351924 pvsat_ff=7.84794e-11                pvsat_ss=-2.35437e-10               pvsat_fs=1.56958e-10 pvsat_sf=-1.56958e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.25 nmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.37587324 lvth0=-1.3200651e-009            wvth0=-9.9501047e-009            pvth0=-2.9337426e-017 k2=-0.02068891                lk2=-1.0886224e-010            wk2=2.722167e-009 pk2=4.3384876e-017             cit=0.0036001527               lcit=-5.526946e-011 wcit=-1.1774347e-010            pcit=1.1371828e-017             voff=-0.1578541 lvoff=-4.5382033e-009            wvoff=1.6433154e-010             pvoff=2.7133852e-016 eta0=0.0036316061               weta0=4.9799691e-010             etab=-0.034056674 wetab=7.1958209e-010             u0=0.019830765                wu0=1.9410991e-010 ua=-1.4860914e-009            lua=-1.5761346e-017            wua=-5.4853445e-017 pua=6.2477797e-024             ub=1.6815347e-018             lub=1.6698839e-026 wub=5.0494423e-026             pub=-6.9904105e-033            uc=7.3565861e-011 wuc=1.9987278e-018             vsat=134595.92                  a0=4.6418894 la0=-6.4722626e-007            wa0=-8.1667116e-008            pa0=4.5506311e-015 ags=2.7857245                  lags=-6.757229e-008             wags=6.3875028e-008 pags=-5.4932541e-015            keta=0.030718141                lketa=-1.9684022e-008 wketa=-7.5099234e-009            pketa=8.3911392e-016             pclm=0.61933702 lpclm=5.2738091e-008             wpclm=3.4512922e-008             ppclm=-1.8290927e-015 pdiblc2=0.0022692014               lpdiblc2=-2.7610576e-011            wpdiblc2=6.0511045e-011 ppdiblc2=3.1476057e-018             aigbacc=0.012884843                laigbacc=5.8307448e-011 waigbacc=-3.5786002e-012            paigbacc=-8.7123864e-018            aigc=0.010666309 laigc=4.520536e-012              waigc=1.8493892e-011             paigc=-5.0489607e-019 aigsd=0.0098181777               laigsd=-1.5075191e-011            waigsd=7.9292264e-012 paigsd=-3.0503783e-019            tvoff=0.00228564                 ltvoff=-1.26937e-010 wtvoff=-1.43705e-010              ptvoff=2.30486e-017               kt1=-0.18191949 lkt1=5.1006635e-009             wkt1=-2.1582352e-009            pkt1=1.1265572e-016 kt2=-0.069501513               lkt2=7.5198642e-010             wkt2=-3.3538236e-010 pkt2=-1.6561465e-016            ute=-1.1127668                 lute=8.3484553e-010 wute=-9.4827983e-009            pute=4.0629443e-016             ua1=1.6253577e-009 lua1=-9.6087631e-017            wua1=-1.0496306e-016            pua1=5.0417952e-024 ub1=-1.489964e-018             lub1=6.9779e-026                wub1=9.7323511e-026 pub1=-4.6763117e-033            uc1=5.5068783e-011             luc1=5.7879365e-018 wuc1=1.5537778e-018             puc1=-1.3066393e-039            at=66886.244 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=-1.4726212e-009            petab=-1.525514e-016             lu0=8.595761e-012 pu0=-3.8627901e-018            luc=-7.3430802e-019            puc=-2.414787e-025 lat=-0.00098902673             wat=0.0051771485               pat=-3.5220413e-010 lvsat=-0.0020186319              wvsat=0.00044625012              pvsat=1.9362075e-010 leta0=6.6871892e-010             peta0=-7.6233956e-017            vsat_ff=-7072.88 vsat_ss=8599.65                    vsat_fs=-5733.1                    vsat_sf=5733.1 a0_ff=1.08312                    a0_ss=-1.5766                    a0_fs=0.914051 a0_sf=-0.859965                  la0_ff=-6.00236e-08               la0_ss=1.35588e-07 la0_fs=-4.93047e-08               la0_sf=7.3957e-08                 wa0_ff=6.62899e-09 wa0_ss=1.79733e-07                wa0_fs=-1.04202e-07               wa0_sf=9.8036e-08 pa0_ff=-1.40523e-15               pa0_ss=-1.5457e-14                pa0_fs=5.62077e-15 pa0_sf=-8.43109e-15               pdiblc2_ff=-5.92005e-05               pdiblc2_fs=5.92005e-05 lpdiblc2_ff=5.09124e-12                lpdiblc2_fs=-5.09124e-12               wpdiblc2_ff=1.63393e-11 wpdiblc2_fs=-1.63393e-11               ppdiblc2_ff=-1.40518e-18               ppdiblc2_fs=1.40518e-18 lvsat_ff=0.000608269                lvsat_ss=-0.00073957                lvsat_fs=0.000493046 lvsat_sf=-0.000493046               wvsat_ff=0.000326784                wvsat_ss=-0.00098036 wvsat_fs=0.000653573                wvsat_sf=-0.000653573               pvsat_ff=-2.81037e-11 pvsat_ss=8.43109e-11                pvsat_fs=-5.62073e-11               pvsat_sf=5.62073e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.26 nmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.35455727 lvth0=5.1310821e-010             wvth0=-1.1565637e-008            pvth0=1.0959832e-016 k2=-0.018938758               lk2=-2.5937531e-010            wk2=2.7908878e-009 pk2=3.7474892e-017             cit=-2.1057646e-005            lcit=2.5615463e-010 wcit=2.4868025e-010             pcit=-2.0140611e-017            voff=-0.20426941 lvoff=-5.4648654e-010            wvoff=5.3855313e-009             pvoff=-1.7768466e-016 eta0=0.0056874538               weta0=1.9712792e-010             etab=-0.074503353 wetab=-2.9691431e-009            u0=0.021831198                wu0=6.9595811e-011 ua=-1.9076976e-009            lua=2.0496792e-017             wua=8.5662642e-018 pua=7.9368475e-025             ub=2.0156916e-018             lub=-1.2038656e-026 wub=-3.1077616e-026            pub=2.4784865e-035             uc=5.1094621e-012 wuc=4.5106424e-018             vsat=85280.601                  a0=-1.4358867 la0=-1.2453751e-007            wa0=8.9292858e-007             pa0=-7.9264599e-014 ags=2.0000004                  lags=-2.0349794e-014            wags=-4.639753e-014 pags=2.3198765e-021             keta=-0.44845696                lketa=2.1525037e-008 wketa=4.0651796e-008             pketa=-3.3027939e-015            pclm=1.2778076 lpclm=-3.8903817e-009            wpclm=3.1639404e-008             ppclm=-1.5819702e-015 pdiblc2=0.0026580247               lpdiblc2=-6.1049383e-011            wpdiblc2=1.6185185e-011 ppdiblc2=6.9596296e-018             aigbacc=0.016469096                laigbacc=-2.4993828e-010 waigbacc=-5.4907428e-010            paigbacc=3.8200242e-017             aigc=0.010878608 laigc=-1.3737145e-011            waigc=1.9310429e-011             paigc=-5.7511827e-019 aigsd=0.0096825095               laigsd=-3.4077266e-012            waigsd=-4.7223612e-012 paigsd=7.829987e-019              tvoff=-0.000884274               ltvoff=1.45676e-010 wtvoff=4.2824e-010                ptvoff=-2.61387e-017              kt1=-0.13678794 lkt1=1.2193497e-009             wkt1=7.6562076e-010             pkt1=-1.3879589e-016 kt2=-0.056161811               lkt2=-3.9522798e-010            wkt2=-3.1270402e-009 pkt2=7.4467921e-017             ute=-1.1773288                 lute=6.3871811e-009 wute=-9.1716049e-011            pute=-4.0133864e-016            ua1=2.7790587e-010 lua1=1.9793224e-017             wua1=-2.1083261e-017            pua1=-2.171868e-024 ub1=-5.2368389e-020            lub1=-5.385422e-026             wub1=-3.1491305e-027 pub1=3.9643354e-033             uc1=1.4911934e-010             luc1=-2.3004115e-018 wuc1=-2.7622716e-018            puc1=3.7118025e-025             at=40113.86 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=2.0057932e-009             petab=1.6467897e-016             lu0=-1.6344142e-010 pu0=6.8454221e-018             luc=5.1529423e-018             puc=-4.5750337e-025 lat=0.0013133983               wat=0.0023472182               pat=-1.0883012e-010 lvsat=0.0022224857               wvsat=0.0053683495               pvsat=-2.296798e-010 leta0=4.9191601e-010             peta0=-5.0359223e-017            vsat_ff=1388.89 a0_ff=0.920169                   a0_fs=0.813992                   la0_ff=-4.60083e-08 la0_fs=-4.06996e-08               wa0_ff=-2.31984e-08               wa0_fs=-9.27951e-08 pa0_ff=1.15994e-15                pa0_fs=4.63975e-15                lvsat_ff=-0.000119445 wvsat_ff=9e-11                      pvsat_ff=3.5e-17 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.27 nmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.444148 lvth0=-3.9664283e-009            wvth0=-1.9213348e-008            pvth0=4.9198388e-016 k2=-0.016321194               lk2=-3.9025352e-010            wk2=2.4827067e-009 pk2=5.2883945e-017             cit=0.00049924727              lcit=2.3013938e-010 wcit=8.1592391e-011             pcit=-1.1786218e-017            voff=-0.28812398 lvoff=3.6462423e-009             wvoff=1.3825923e-008             pvoff=-5.9970424e-016 eta0=-0.0084941693              weta0=-2.2679887e-009            etab=-0.076849927 wetab=-1.0121246e-010            u0=0.019124355                wu0=3.7410828e-010 ua=-2.4858226e-009            lua=4.9403041e-017             wua=1.1073941e-016 pua=-4.3149723e-024            ub=2.0629055e-018             lub=-1.439935e-026 wub=-3.3496815e-026            pub=1.4574484e-034             uc=1.0182785e-010 wuc=1.3336694e-018             vsat=190901.68                  a0=12.677964 la0=-8.3023002e-007            wa0=-2.7054716e-006            pa0=1.0065541e-013 ags=2                          lags=0                          wags=0 pags=0                          keta=0.14009556                 lketa=-7.9025889e-009 wketa=-6.9026374e-008            pketa=2.1811145e-015             pclm=0.87942387 lpclm=1.6028807e-008             wpclm=8.8479012e-008             ppclm=-4.4239506e-015 pdiblc2=0.001437037                lpdiblc2=0                          wpdiblc2=1.5537778e-010 ppdiblc2=0                          aigbacc=0.001358751                laigbacc=5.0557897e-010 waigbacc=1.8120289e-009             paigbacc=-7.9854919e-017            aigc=0.010656976 laigc=-2.655554e-012             waigc=1.1592222e-011             paigc=-1.8920794e-019 aigsd=0.0091004108               laigsd=2.5697209e-011             waigsd=8.2720034e-011 paigsd=-3.5891211e-018            tvoff=0.00580062                 ltvoff=-1.88569e-010 wtvoff=-6.95849e-010              ptvoff=3.00658e-017               kt1=0.10476852 lkt1=-1.0858473e-008            wkt1=-2.6635565e-008            pkt1=1.2312634e-015 kt2=-0.14944846                lkt2=4.2691043e-009             wkt2=8.7284229e-009 pkt2=-5.1830523e-016            ute=-0.76442259                lute=-1.425813e-008 wute=-4.2773948e-008            pute=1.732773e-015              ua1=8.2654654e-010 lua1=-7.6388089e-018            wua1=-1.8212687e-016            pua1=5.8803125e-024 ub1=-6.9333433e-019            lub1=-2.1805924e-026            wub1=1.724968e-025 pub1=-4.8179609e-033            uc1=4.3920988e-010             luc1=-1.6804938e-017 wuc1=-3.7808593e-017            puc1=2.1234963e-024             at=54227.15 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=2.1231219e-009             petab=2.1282432e-017             lu0=-2.8099308e-011 pu0=-8.3802012e-018            luc=3.1702275e-019             puc=-2.9865471e-025 lat=0.00060773384              wat=-0.0062968723              pat=3.2337441e-010 lvsat=-0.0030585684              wvsat=-0.014314391               pvsat=7.5445722e-010 leta0=1.2009972e-009             peta0=7.2896605e-017             uc_ss=-9.61728e-11 wuc_ss=2.65437e-17                vsat_ff=-5555.56                   vsat_fs=-7761.32 ua1_ss=-2.24403e-10               lua1_ss=1.12202e-17                wua1_ss=6.19353e-17 pua1_ss=-3.09677e-24               uc1_sf=2.88519e-10                uc1_ss=4.80864e-10 luc1_sf=-1.44259e-17               luc1_ss=-2.40432e-17               wuc1_sf=-7.96311e-17 wuc1_ss=-1.32719e-16               puc1_sf=3.98156e-24                puc1_ss=6.63593e-24 luc_ss=4.80864e-18                puc_ss=-1.32719e-24               lvsat_ff=0.000227778 lvsat_fs=0.000388066                wvsat_ff=-2.3e-09                   wvsat_fs=0.00088479 pvsat_ff=6e-18                      pvsat_fs=-4.42395e-11 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_lvt_mac.28 nmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=0.33797475 lvth0=3.8667493e-010             wvth0=-1.0630516e-008            pvth0=1.4008779e-016 k2=0.0092585175               lk2=-1.4390217e-009            wk2=2.87052e-009 pk2=3.69836e-017               cit=-0.015373998               lcit=8.8094243e-010 wcit=1.1773372e-009             pcit=-5.6711754e-017            voff=-0.048327923 lvoff=-6.1853962e-009            wvoff=-1.2208428e-008            pvoff=4.6770417e-016 eta0=-0.0058674321              weta0=1.0906873e-009             etab=-0.052943508 wetab=9.2380961e-010             u0=0.018908485                wu0=2.5039148e-010 ua=-1.3534761e-009            lua=2.9768372e-018             wua=-4.3415745e-017 pua=2.0053889e-024             ub=1.8320815e-018             lub=-4.9355663e-027 wub=-7.2344226e-027            pub=-9.3101326e-034            uc=2.8578932e-010 wuc=-9.6634102e-018            vsat=-13615.348                 a0=0.49340604 la0=-3.3066316e-007            wa0=-1.0760645e-006            pa0=3.3849719e-014 ags=2                          lags=0                          wags=0 pags=0                          keta=-0.050096327               lketa=-1.0472168e-010 wketa=-5.9425819e-008            pketa=1.7874918e-015             pclm=3.4958848 lpclm=-9.124609e-008             wpclm=-1.920642e-007             ppclm=7.0783213e-015 pdiblc2=0.001437037                lpdiblc2=0                          wpdiblc2=1.5537778e-010 ppdiblc2=0                          aigbacc=0.015537786                laigbacc=-7.5761474e-011 waigbacc=-2.2963816e-010            paigbacc=3.8534323e-018             aigc=0.010514911 laigc=3.1691106e-012             waigc=7.0396872e-011             paigc=-2.6001986e-018 aigsd=0.010034351                laigsd=-1.2594356e-011            waigsd=-9.0214268e-011 paigsd=3.5011853e-018             tvoff=0.00268797                 ltvoff=-6.09502e-011 wtvoff=6.59561e-011               ptvoff=-1.16824e-018              kt1=-0.054860391 lkt1=-4.3136879e-009            wkt1=-2.6362105e-009            pkt1=2.4728986e-016 kt2=0.0068575163               lkt2=-2.1394406e-009            wkt2=-1.7826657e-008 pkt2=5.7045304e-016             ute=-0.96737988                lute=-5.936881e-009 wute=-1.6761637e-008            pute=6.662682e-016              ua1=5.0616382e-010 lua1=5.4968827e-018             wua1=-4.7727724e-018            pua1=-1.3912055e-024 ub1=-2.0149413e-018            lub1=3.2379964e-026             wub1=1.6642548e-025 pub1=-4.5690369e-033            uc1=-2.3614815e-010            luc1=1.0884741e-017 wuc1=6.3704889e-017             puc1=-2.0385564e-024            at=-67026.485 jtsswgs='5.2e-006*(1+1.55*iboffn_flag_lvt)'                                jtsswgd='5.2e-006*(1+1.55*iboffn_flag_lvt)' letab=1.1429587e-009             petab=-2.0743473e-017            lu0=-1.9248644e-011 pu0=-3.3078126e-018            luc=-7.2253972e-018            puc=1.5222555e-025 lat=0.0055791328               wat=0.012810779                pat=-4.6003931e-010 lvsat=0.0053266299               wvsat=0.010203884                pvsat=-2.5079205e-010 leta0=1.0933009e-009             peta0=-6.4809107e-017            cit_mcl=-0.00605761 lcit_mcl=2.48362e-10                wcit_mcl=6.90568e-10                pcit_mcl=-2.83133e-17 voff_ff=-0.0302881                 lvoff_ff=1.24181e-09                wvoff_ff=3.45284e-09 pvoff_ff=-1.41566e-16               u0_ss=-0.00363457                u0_ff=0.00212016 u0_sf=-0.00121152                wu0_ss=4.14341e-10                wu0_ff=-2.41699e-10 wu0_sf=1.38114e-10                uc_ss=9.61728e-11                wuc_ss=-2.65437e-17 vsat_ss=-18172.8                   vsat_ff=24230.5                    vsat_sf=-12115.2 vsat_fs=7761.32                    ua1_ss=2.24403e-10                lua1_ss=-7.18091e-18 wua1_ss=-6.19353e-17               pua1_ss=1.98193e-24                uc1_sf=-3.63581e-10 uc1_ss=-5.80946e-10               luc1_sf=1.23101e-17                luc1_ss=1.94911e-17 wuc1_sf=1.00348e-16                wuc1_ss=1.60342e-16                puc1_sf=-3.3976e-24 puc1_ss=-5.37952e-24               lu0_ss=1.49017e-10                lu0_ff=-8.69267e-11 lu0_sf=4.96724e-11                pu0_ss=-1.6988e-17                pu0_ff=9.90965e-18 pu0_sf=-5.66266e-18               luc_ss=-3.07753e-18               puc_ss=8.49399e-25 lvsat_ss=0.000745086                lvsat_ff=-0.000993449               lvsat_sf=0.000496724 lvsat_fs=-0.000248362               wvsat_ss=0.0020717                  wvsat_ff=-0.00276227 wvsat_sf=0.00138114                 wvsat_fs=-0.00088479                pvsat_ss=-8.49399e-11 pvsat_ff=1.13253e-10                pvsat_sf=-5.66266e-11               pvsat_fs=2.83133e-11 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model pch_lvt_mac.global pmos ( modelid=6                          level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_lvt'             permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          wpemod=1 tnom=25                         toxe=2.18e-009                  toxm=2.18e-009 dtox=4.422e-010                 epsrox=3.9                        toxref=3e-009 wint=0                          lint=0                          ll=0 wl=0                          lln=1                          wln=1 lw=0                          ww=0                          lwn=1 wwn=1                          lwl=0                          wwl=0 llc=0                          wlc=0                          lwc=0 wwc=0                          lwlc=0                          wwlc=0 xl=-3e-009                    xw=6e-009                     dlc=7.64e-009 dwc=0                          dlcig=2.5e-009                   xpart=1 k1=0.34                       k3=-2.45                      k3b=2.25 w0=0                          dvt0=20                         dvt1=2.5853 dvt2=-0.14                      dvt0w=0                          dvt1w=0 dvt2w=0                          dsub=0.5                        minv=-0.3292 voffl=0                          dvtp0=1.478e-007                 dvtp1=0.3 lpe0=1e-010                     lpeb=-2.5e-008                  xj=8.5e-008 ngate=1.17e+020                  ndep=6e+017                     nsd=1e+020 phin=0.15                       cdsc=0                          ud=0 cdscb=0                          cdscd=0                          nfactor=0.8 a1=0                          a2=1                          b0=0 b1=0                          dwg=0                          dwb=0 pdiblc1=0                          pdiblcb=0                          drout=0.56 pvag=0.07                       delta=0.015992                   pscbe1=9.264e+008 pscbe2=1e-020                     fprout=200                        pdits=0 pditsd=0                          pditsl=0                          rsh=16.7 rdsw=160                        prwg=0                          prwb=0 wr=1                          alpha0=1.5675e-006                alpha1=2 beta0=18.727                     agidl=1e-008                     bgidl=2.2565e+009 cgidl=8                          egidl=0.001                      bigbacc=0.006 cigbacc=0.245                      nigbacc=10                         aigbinv=0.009974 bigbinv=0.00149                    cigbinv=0.006                      eigbinv=1.1 nigbinv=2.171                      bigc=0.0013746                  cigc=0.15259 bigsd=0.00024                    cigsd=0.0011                     nigc=2.291 poxedge=1                          pigcd=3                          ntox=1 vfbsdoff=0.01                       cgso=5.71e-011                  cgdo=5.71e-011 cgbo=0                          cgdl=6.7e-011                   cgsl=6.7e-011 clc=0                          cle=0.6                        cf='9e-011+9.2e-11*ccoflag_lvt' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=6                          noff=2.4                        voffcv=-0.1 tvfbsdoff=0.114                      kt1l=0                          prt=0 fnoimod=1                          tnoimod=0                          em=5.63e+006 ef=1.12                       noia=0                          noib=0 noic=0                          lintnoi=-3.26e-008                 jss=3.97e-07 jsd=3.97e-07                   jsws=8.37e-14                   jswd=8.37e-14 jswgs=8.37e-14                   jswgd=8.37e-14                   njs=1.02 njd=1.02                       ijthsfwd=0.01                       ijthdfwd=0.01 ijthsrev=0.01                       ijthdrev=0.01                       bvs=7.58 bvd=7.58                       xjbvs=1                          xjbvd=1 njtsswg=36                         xtsswgs=0.1                        xtsswgd=0.1 tnjtsswg=1                          vtsswgs=1                          vtsswgd=1 pbs=0.778                      pbd=0.778                      cjs=0.001474 cjd=0.001474                   mjs=0.421                      mjd=0.421 pbsws=0.751                      pbswd=0.751                      cjsws=1.07e-010 cjswd=1.07e-010                  mjsws=0.254                      mjswd=0.254 pbswgs=0.944                      pbswgd=0.944                      cjswgs=2.07e-010 cjswgd=2.07e-010                  mjswgs=0.672                      mjswgd=0.672 tpb=0.00104                    tcj=0.00079                    tpbsw=0.00089 tcjsw=0.00030                    tpbswg=0.00214                    tcjswg=0.00170 xtis=3                          xtid=3                          dmcg=3.75e-008 dmci=3.75e-008                  dmdg=0                          dmcgt=0 dwj=0                          xgw=0                          xgl=-5.1e-009 rshg=14.4                       gbmin=1e-012                     rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         ngcon=1                          xrcrg1=12 xrcrg2=1                          web=2251.7                     wec=-7896.1 scref=1e-6                       kvth0we=-0.0004346                 k2we=0.0000 ku0we=-0.0007                    lk2we=0                          lku0we=-2e-11 lkvth0we=10e-012                    pk2we=0                          pku0we=4.5e-18 pkvth0we=0e-019                     wk2we=0                          wku0we=-1.3e-10 wkvth0we=-1e-011 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.1                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.2                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.1 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.6 bidirectionflag='bidirectionflag_mos_lvt' iboffn_flag='iboffn_flag_lvt' iboffp_flag='iboffp_flag_lvt' sigma_factor='sigma_factor_lvt' ccoflag='ccoflag_lvt' rcoflag='rcoflag_lvt' rgflag='rgflag_lvt' mismatchflag='mismatchflag_mos_lvt' globalflag='globalflag_mos_lvt' totalflag='totalflag_mos_lvt' designflag='designflag_mos_lvt' global_factor='global_factor_lvt' local_factor='local_factor_lvt' sigma_factor_flicker='sigma_factor_flicker_lvt' noiseflag='noiseflagp_lvt' noiseflag_mc='noiseflagp_lvt_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w51='2.3875*0.35355' w52='0.70711*0.35355' w53='0.54772*0.22143' w54='0.54772*-0.066279' w55='0.54772*0.050463' w56='0.54772*-0.03945' w57='0.54772*-0.80208' w58='0.54772*0.22166' w59='0' w60='0' tox_c='toxp_lvt'                 dxl_c='dxlp_lvt'                 dxw_c='dxwp_lvt' cgo_c='cgop_lvt'                 cgl_c='cglp_lvt'                 ddlc_c='ddlcp_lvt' cj_c='cjp_lvt'                  cjsw_c='cjswp_lvt'                cjswg_c='cjswgp_lvt' cf_c='cfp_lvt'                  dvth_c='dvthp_lvt'                dlvth_c='dlvthp_lvt' dwvth_c='dwvthp_lvt'               dpvth_c='dpvthp_lvt'               dk2_c='dk2p_lvt' dlk2_c='dlk2p_lvt'                dwk2_c='dwk2p_lvt'                dpk2_c='dpk2p_lvt' deta0_c='deta0p_lvt'               dweta0_c='dweta0p_lvt'              dvoff_c='dvoffp_lvt' dlvoff_c='dlvoffp_lvt'              dwvoff_c='dwvoffp_lvt'              dpvoff_c='dpvoffp_lvt' du0_c='du0p_lvt'                 dlu0_c='dlu0p_lvt'                dwu0_c='dwu0p_lvt' dpu0_c='dpu0p_lvt'                dpclm_c='dpclmp_lvt'               dlpclm_c='dlpclmp_lvt' dwpclm_c='dwpclmp_lvt'              dppclm_c='dppclmp_lvt'              dpdiblc2_c='dpdiblc2p_lvt' dwpdiblc2_c='dwpdiblc2p_lvt'           dlpdiblc2_c='dlpdiblc2p_lvt'           dppdiblc2_c='dppdiblc2p_lvt' da0_c='da0p_lvt'                 dla0_c='dla0p_lvt'                dwa0_c='dwa0p_lvt' dpa0_c='dpa0p_lvt'                dags_c='dagsp_lvt'                dlags_c='dlagsp_lvt' dwags_c='dwagsp_lvt'               dpags_c='dpagsp_lvt'               ntox_c='ntoxp_lvt' dvsat_c='dvsatp_lvt'               dlvsat_c='dlvsatp_lvt'              dwvsat_c='dwvsatp_lvt' dpvsat_c='dpvsatp_lvt'              dminv_c='dminvp_lvt'               dat_c='datp_lvt' dua1_c='dua1p_lvt'                dlua1_c='dlua1p_lvt'               dwua1_c='dwua1p_lvt' dpua1_c='dpua1p_lvt'               jtsswg_c='jtsswgp_lvt'              ss_flag_c='ss_flagp_lvt' ff_flag_c='ff_flagp_lvt'             sf_flag_c='sf_flagp_lvt'             fs_flag_c='fs_flagp_lvt' monte_flag_c='monte_flagp_lvt'         c1f_c='c1fp_lvt'                 c2f_c='c2fp_lvt' c3f_c='c3fp_lvt' global_mc='global_mc_flag_lvt' tox_g='toxp_lvt_ms_global'       dxl_g='dxlp_lvt_ms_global'       dxw_g='dxwp_lvt_ms_global' cgo_g='cgop_lvt_ms_global'       cgl_g='cglp_lvt_ms_global'       cj_g='cjp_lvt_ms_global' cjsw_g='cjswp_lvt_ms_global'      cjswg_g='cjswgp_lvt_ms_global'     cf_g='cfp_lvt_ms_global' dvth_g='dvthp_lvt_ms_global'      dlvth_g='dlvthp_lvt_ms_global' dwvth_g='dwvthp_lvt_ms_global'     dpvth_g='dpvthp_lvt_ms_global'     dk2_g='dk2p_lvt_ms_global' dlk2_g='dlk2p_lvt_ms_global'      dwk2_g='dwk2p_lvt_ms_global'      dpk2_g='dpk2p_lvt_ms_global' deta0_g='deta0p_lvt_ms_global'     dvoff_g='dvoffp_lvt_ms_global' dlvoff_g='dlvoffp_lvt_ms_global'    du0_g='du0p_lvt_ms_global'       dlu0_g='dlu0p_lvt_ms_global' dwu0_g='dwu0p_lvt_ms_global'      dpu0_g='dpu0p_lvt_ms_global' dpclm_g='dpclmp_lvt_ms_global'     dpdiblc2_g='dpdiblc2p_lvt_ms_global' dags_g='dagsp_lvt_ms_global'      dwags_g='dwagsp_lvt_ms_global' ntox_g='ntoxp_lvt_ms_global'      dvsat_g='dvsatp_lvt_ms_global' dlvsat_g='dlvsatp_lvt_ms_global'    dwvsat_g='dwvsatp_lvt_ms_global' dpvsat_g='dpvsatp_lvt_ms_global'    dminv_g='dminvp_lvt_ms_global'     dat_g='datp_lvt_ms_global' dua1_g='dua1p_lvt_ms_global'      dlua1_g='dlua1p_lvt_ms_global' ss_flag_g='ss_flagp_lvt_ms_global'   ff_flag_g='ff_flagp_lvt_ms_global' monte_flag_g='monte_flagp_lvt_ms_global'                                       sf_flag_g='sf_flagp_lvt_ms_global' fs_flag_g='fs_flagp_lvt_ms_global' weight1=-3.2374522 weight2=2.0282803 weight3=-0.98369427 weight4=0.63694268 weight5=-0.44434395 tox_1=4.3392818e-012 tox_2=-9.4753602e-012 tox_3=-9.6435595e-013 tox_4=-3.7476843e-011 tox_5=5.4457771e-013 dxl_1=9.8246587e-011 dxl_2=-2.145391e-010 dxl_3=-2.1834908e-011 dxl_4=8.4852644e-010 dxl_5=1.2329948e-011 dxl_max=-2e-009 dxw_1=-6.8725711e-010 dxw_2=-8.2201655e-010 dxw_3=6.186374e-011 dxw_4=5.1808782e-025 dxw_5=-5.8973752e-009 cgo_1=-3.8811e-013 cgo_2=9.6993e-014 cgo_3=5.265e-014 cgo_4=1.2149e-028 cgo_5=3.3278e-014 cgl_1=-4.554e-013 cgl_2=1.1381e-013 cgl_3=6.1779e-014 cgl_4=7.2035e-029 cgl_5=3.9048e-014 cj_1=1.0019e-005 cj_2=-2.5038e-006 cj_3=-1.3591e-006 cj_4=9.6855e-022 cj_5=-8.5905e-007 cjsw_1=7.2727e-013 cjsw_2=-1.8176e-013 cjsw_3=-9.8661e-014 cjsw_4=-3.7803e-028 cjsw_5=-6.236e-014 cjswg_1=1.407e-012 cjswg_2=-3.5162e-013 cjswg_3=-1.9087e-013 cjswg_4=-7.3132e-028 cjswg_5=-1.2064e-013 cf_1=-6.1173e-013 cf_2=1.5288e-013 cf_3=8.2986e-014 cf_4=-7.2245e-029 cf_5=5.2452e-014 dvth_1=-0.0032965 dvth_2=-0.0026592 dvth_3=0.00029125 dvth_4=1.2104e-018 dvth_5=0.00066316 dlvth_1=-9.1444e-011 dlvth_2=-8.1851e-011 dlvth_3=2.286e-011 dlvth_4=-1.188e-025 dlvth_5=1.9884e-011 dwvth_1=-1.4037e-010 dwvth_2=1.7162e-011 dwvth_3=3.6191e-011 dwvth_4=3.1867e-026 dwvth_5=1.2988e-011 dpvth_1=-2.4174e-017 dpvth_2=-9.8036e-018 dpvth_3=4.4274e-018 dpvth_4=-8.2198e-033 dpvth_5=3.819e-018 dk2_1=0.00015943 dk2_2=-4.3808e-005 dk2_3=0.00054257 dk2_4=2.9679e-019 dk2_5=-8.5988e-006 dlk2_1=9.0493e-012 dlk2_2=-2.421e-012 dlk2_3=2.1483e-011 dlk2_4=-3.3742e-027 dlk2_5=-5.7177e-013 dwk2_1=1.4195e-010 dwk2_2=-3.6177e-011 dwk2_3=8.0728e-011 dwk2_4=7.0598e-026 dwk2_5=-1.1272e-011 dpk2_1=-1.8874e-018 dpk2_2=4.8283e-019 dpk2_3=-1.3294e-018 dpk2_4=-7.134e-035 dpk2_5=1.4759e-019 deta0_1=-0.00097099 deta0_2=0.00024266 deta0_3=0.00013172 deta0_4=-3.4706e-019 deta0_5=8.3258e-005 dvoff_1=-0.0004855 dvoff_2=0.00012133 dvoff_3=6.5862e-005 dvoff_4=-2.9109e-019 dvoff_5=4.1629e-005 dlvoff_1=7.7679e-011 dlvoff_2=-1.9413e-011 dlvoff_3=-1.0538e-011 dlvoff_4=8.7537e-027 dlvoff_5=-6.6606e-012 du0_1=8.7121e-005 du0_2=9.8812e-005 du0_3=1.7308e-005 du0_4=6.2186e-020 du0_5=-2.2369e-005 dlu0_1=1.6767e-012 dlu0_2=1.0891e-011 dlu0_3=-1.6594e-012 dlu0_4=-3.2866e-027 dlu0_5=-2.3557e-012 dwu0_1=8.1434e-012 dwu0_2=1.2773e-011 dwu0_3=9.285e-013 dwu0_4=1.4052e-026 dwu0_5=-2.0166e-012 dpu0_1=3.1064e-019 dpu0_2=2.912976e-018 dpu0_3=6.6559e-020 dpu0_4=8.0181e-034 dpu0_5=-7.6496e-019 dpclm_1=-0.004855 dpclm_2=0.0012133 dpclm_3=0.00065862 dpclm_4=-2.1234e-018 dpclm_5=0.00041629 dpclm_max=-0.01 dpdiblc2_1=-2.913e-005 dpdiblc2_2=7.2799e-006 dpdiblc2_3=3.9517e-006 dpdiblc2_4=-1.9931e-020 dpdiblc2_5=2.4977e-006 dags_1=0.034138 dags_2=0.027852 dags_3=0.0012844 dags_4=-2.5313e-017 dags_5=-0.0068665 dwags_1=1.8857e-010 dwags_2=1.9228e-009 dwags_3=1.1331e-011 dwags_4=-1.0613e-025 dwags_5=-2.6061e-010 ntox_1=0.01942 ntox_2=-0.0048533 ntox_3=-0.0026345 ntox_4=8.4936e-018 ntox_5=-0.0016652 dvsat_1=212.77 dvsat_2=2174.6 dvsat_3=-14.603 dvsat_4=-8.5697e-013 dvsat_5=-310.34 dlvsat_1=1.1824e-005 dlvsat_2=-3.4509e-005 dlvsat_3=-1.8734e-005 dlvsat_4=-2.2067e-020 dlvsat_5=2.304e-006 dwvsat_1=1.5227e-005 dwvsat_2=0.00015451 dwvsat_3=5.0231e-006 dwvsat_4=4.7446e-021 dwvsat_5=-1.8601e-005 dwvsat_max=0 dpvsat_1=3.3232e-012 dpvsat_2=1.5244e-011 dpvsat_3=-3.7555e-012 dpvsat_4=4.8397e-027 dpvsat_5=-3.0345e-012 dminv_1=-0.011216 dminv_2=0.0028331 dminv_3=-0.0027635 dminv_4=2.5891e-018 dminv_5=0.00092318 dat_1=1456.5 dat_2=-364 dat_3=-197.59 dat_4=1.4297e-012 dat_5=-124.89 dua1_1=2.913e-012 dua1_2=-7.2799e-013 dua1_3=-3.9517e-013 dua1_4=-4.4228e-027 dua1_5=-2.4977e-013 dlua1_1=-1.8761e-019 dlua1_2=4.2874e-020 dlua1_3=5.9679e-019 dlua1_4=2.1158e-034 dlua1_5=2.1223e-020 ss_flag_1=0.050196 ss_flag_2=-0.013548 ss_flag_3=0.13603 ss_flag_4=-1.4407e-016 ss_flag_5=-0.00302 ff_flag_1=-0.046903 ff_flag_2=0.010718 ff_flag_3=0.1492 ff_flag_4=1.1615e-016 ff_flag_5=0.0053057 monte_flag_1=0.0818725 monte_flag_2=-0.178783 monte_flag_3=-0.0181958 monte_flag_4=0.707108 monte_flag_5=0.010275 sigma_local=1                          a_1=0.907705 b_1=-0.00021893                c_1=0.00344948                 d_1=0.00012579 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1.06704                    b_2=-0.00445013                c_2=-0.00712538 d_2=-0.000413874               a_3=0.972014                   b_3=-0.0065125 c_3=-0.00516675                d_3=-0.000203729               e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=1 b_4=-0.0043                    c_4=-0.0015                    d_4=-0.0002 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=0.97                       b_5=-7.5e-3                    c_5=-0.0015 d_5=-0.0002                    e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=-0.00145                   mis_a_2=-0.05                      mis_a_3=0.0 mis_b_1=0.00365                    mis_b_2=0.03                       mis_b_3=0.08 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.0007                     mis_d_2=0                          mis_d_3=0 mis_e_1=0.003                      mis_e_2=0.5                        mis_e_3=0.02 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-3e-09 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=60                         co_rsd=16.7 cf0=9e-011                     cco=9.2e-11 lres=1e-6                       lrdr1=3.6e-008                   lrdr2=4.05e-008 lrdr3=4.5e-008                   lrdr4=5.4e-008                   lrdr5=6.3e-008 lrdr6=7.2e-008                   lrdr_low=7.2e-008                   lrdr_high=9.0009e-006 r_rjtsswg=0.6                        l_rjtsswg=0                          ll_rjtsswg=0.0 w_rjtsswg=5.0e-04                    ww_rjtsswg=3.0                        p_rjtsswg=0.0 noimod=1                          noic2='2.236'                    noic3='0.5' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.261e-6            sbref0=0.261e-6 samax=10e-6               sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=1                   lreflod=0.9e-6              llodref=2 lod_clamp=-1e90 wlod0=0 ku00=-0e-9       lku00=0e-7        wku00=0e-8         pku00=0e-14 tku00=0           llodku00=1           wlodku00=1            kvsat0=0.5 kvth00=-3.8e-9     lkvth00=1.75e-8     wkvth00=3e-8         pkvth00=0e-15 llodvth0=1           wlodvth0=1 stk20=0           lodk20=1           steta00=5e-11        lodeta00=1 wlod00=0 ku000=0           lku000=-13e-32     wku000=0            pku000=0 llodku000=3           wlodku000=1 kvth000=0           lkvth000=3e-17       wkvth000=0            pkvth000=0e-14 llodvth00=1           wlodvth00=1 steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0           llod1=0.00e-6 ku01=2e-8        lku01=-3e-2       wku01=-5e-15     pku01=0 llodku01=-1          wlodku01=1           kvsat1=-0 kvth01=11e-9     lkvth01=-3e-24      wkvth01='1.5e-19'     pkvth01=0e-24 llodvth1=2           wlodvth1=1.5 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.1        lku02=0.4e-7      wku02=0            pku02=0 tku02=0           llodku02=1           wlodku02=1            kvsat2='0.4*0+0.5' kvth02=-0e-3       lkvth02=0e-8        wkvth02=0e-8         pkvth02=0 llodvth2=1           wlodvth2=1 stk22=0           lodk22=1           steta02=-1e-4        lodeta02=1 wlod02=0 ku002=0           lku002='-1.2e11*2'     wku002=3.5e-9       pku002=0 llodku002=-2          wlodku002=1 kvth002=0           lkvth002=-0e-11      wkvth002=0            pkvth002=0 llodvth02=1           wlodvth02=1 steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0.085        lku03=-0.05e-7        wku03=0e-7         pku03=0 tku03=0           llodku03=1           wlodku03=1            kvsat3=0.4 kvth03=0.1e-3      lkvth03=0e-20       wkvth03=0e-8         pkvth03=0e-20 llodvth3=3           wlodvth3=1 stk23=0           lodk23=1           steta03=0e-3         lodeta03=1 wlod03=0 ku003=0           lku003='-1.25e5*8e-1'     wku003=1.5e-9            pku003=0 llodku003=-1          wlodku003=1 kvth003=0e-3        lkvth003=-5e-26      wkvth003=-2e-10       pkvth003=0e-32 llodvth03=3           wlodvth03=1 steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=2.61e-7             sa_b1=0.99e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.26e-7             spamax=2.88e-7             spamin=1.08e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.7                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=-1.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=-0.000              wkvth0dpl=0                   wdplkvth0=1 lkvth0dpl=0.0e-9              ldplkvth0=1.0                 pkvth0dpl=0 ku0dpl=1               wku0dpl=0                   wdplku0=1 lku0dpl=-4e-8              ldplku0=1                 pku0dpl=0 keta0dpl=0.00                wketa0dpl=0                   wdplketa0=1 kvsatdpl=0                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=1 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=1.0e-6              wkvth0dpx=0                   wdpxkvth0=1 lkvth0dpx=0                   ldpxkvth0=1                   pkvth0dpx=0 ku0dpx=0                   wku0dpx=0                   wdpxku0=1 lku0dpx=0                   ldpxku0=1                   pku0dpx=0 keta0dpx=0                   wketa0dpx=0                   wdpxketa0=1 kvsatdpx=0                   wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0.02               wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-2             ldpskvth0=1.0                 pkvth0dps=0 ku0dps='0.5'               wku0dps=0                   wdpsku0=1 lku0dps='2e-8+0e-8'        ldpsku0=1.0                 pku0dps=0 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0.7                 wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=1 ku0dps_b1=0                 ku0dps_b2=0.11 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=0.002               wkvth0dpa=-2.0e-9            wdpakvth0=1 lkvth0dpa=0.015e-7            ldpakvth0=1.0                pkvth0dpa=-3.0e-17 ku0dpa=-0.1               wku0dpa=2e-9               wdpaku0=1 lku0dpa=-7e-9               ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0                   wka0dpa=0                   wdpaka0=1 lka0dpa=0                   ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=1 ku0dpa_b1=-0.1             ku0dpa_b2=0.00 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=2.88e-7             spbmax='2.88e-7+3.24e-7'    spbmin='1.08e-7+1.38e-7' pse_mode=1 kvth0dp2=-0.01               wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0.5e-9              ldp2kvth0=1                   pkvth0dp2=0 ku0dp2=0.1                wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=-0.0e-8              ldp2ku0=1.0                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0.00                wdp2=0 kvth0dp2l=-0.018              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.6               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0e-8               ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0.2                wdp2l=0 kvth0dp2l_b1=0.00            kvth0dp2l_b2=-0.016           dp2lbinflg=1 ku0dp2l_b1=-0.00            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=-0.007              wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=-0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.2              wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=-25.0e-5            ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=0.017           kvth0dp2a_b2=-0.02           dp2abinflg=1 ku0dp2a_b1=-0.12                ku0dp2a_b2=0.08 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1.44e-7 kvth0enx=-0.023              wkvth0enx=-0.0e-9             wenxkvth0=1.0 lkvth0enx=-11.0e-9              lenxkvth0=1.0                 pkvth0enx=-0.85e-16 ku0enx=-2.0                wku0enx=-1.0e-8             wenxku0=1.0 lku0enx=0.4e-7              lenxku0=1.0                 pku0enx=-7.0e-16 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=1.0                 wka0enx=0                   wenxka0=1 lka0enx=0.0e-7              lenxka0=1.0                 pka0enx=0.0e-14 kvsatenx=0.5                 wenx=0                   ku0enx0=-0.20 eny0=0.08e-6 enyref=0.08e-6             enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0.010               wkvth0eny=5.0e-10             wenykvth0=1 lkvth0eny=1.0e-8              lenykvth0=1.0                 pkvth0eny=0 ku0eny=14.0                wku0eny=1.0e-8              wenyku0=1 ku0eny0=0.04                wku0eny0=-1.0e-7             weny0ku0=1 lku0eny=8.0e-6              lenyku0=1.0                 pku0eny=2.0e-16 keta0eny=0e-4                wketa0eny=0                   wenyketa0=1 ka0eny=-0.00               wka0eny=-0.0e-7             wenyka0=1 lka0eny=-0.0e-7             lenyka0=1.0                 pka0eny=-0.0e-14 kvsateny=0.8                 weny=0 kvth0eny1=-6e-4              wkvth0eny1=0.0e-9             weny1kvth0=1 lkvth0eny1=0.0e-6             leny1kvth0=1.0                pkvth0eny1=3.0e-18 ku0eny1=-1.5e-3            wku0eny1=-1.0e-10           weny1ku0=1 lku0eny1=-0.6e-8            leny1ku0=1.0                pku0eny1=-5.5e-17 keta0eny1=0.00               wketa0eny1=0                  weny1keta0=1 ka0eny1=-0.00              wka0eny1=1.0e-8             weny1ka0=1 lka0eny1=4.0e-9             leny1ka0=1.0                pka0eny1=3.0e-15 kvsateny1=-0.0               weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.9027e-5           ringxmin=0.117e-6 kvth0rx=0.045               wkvth0rx=0.0e-6              wrxkvth0=1.0 lkvth0rx=1.0e-9              lrxkvth0=1.0                 pkvth0rx=0e-15 ku0rx=0.05                wku0rx=0.0e-4              wrxku0=1.0 lku0rx=0.0e-7              lrxku0=1.0                 pku0rx=0.0e-14 keta0rx=0.00                wketa0rx=0                   wrxketa0=1 kvsatrx=0.4                 wrx=0                   ku0rx0=0.35 ry_mode=0 ryref=1.8027e-5           ringymax=1.8047e-5           ringymin=0.117e-6 kvth0ry=-0.0025             wkvth0ry=-0.0e-5             wrykvth0=1.0 lkvth0ry='1.0e-8*0'           lrykvth0=1.0                 pkvth0ry=0.0e-16 ku0ry=-0.8                 wku0ry=-0.5e-8             wryku0=1.0 lku0ry=4.0e-7               lryku0=1.0                 pku0ry=-2.0e-16 keta0ry=0.00                 wketa0ry=0                   wryketa0=1 kvsatry=0.7                 wry=0 kvth0ry0='-0.01*0'            ku0ry0='-0.14*0' sfxref=9.0e-8            sfxmax=1.53e-6          minwodx=0 sfxmin=0.072e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=0.0 kvth0odx1a=-0.009            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.07              lku0odx1a=1.6e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.6 kvth0odx1b=0.0000            lkvth0odx1b=2.7e-11           lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=0.0011            lku0odx1b=1.1e-6            lodx1bku0=0.5 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6 sfymax=1.53e-6           minwody=0.0e-6            wody=5e-7 kvth0odya=40                lkvth0odya=1.0e-4            lodyakvth0=1.0 wkvth0odya=1.8e-7            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=1                 lku0odya=1.0e-6            lodyaku0=1.0 wku0odya=-0.0e-8           wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=-1.5e-2           wketa0ody=0                 wodyketa0=1 kvsatody=0.0 lrefody=1.0e-7            lodyref=1 kvth0odyb=-0.00             lkvth0odyb=7.0e-17           lodybkvth0=2.0 wkvth0odyb=9.0e-9            wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.50             lku0odyb=0.6e-10           lodybku0=1.2 wku0odyb=-0.9e-7           wodybku0=1.0               pku0odyb=-1.8e-16 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=1 oseflag=1 wpeflag=1 )
.model pch_lvt_mac.1 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.34715453 lvth0=-3.3181741e-008            wvth0=-4.211654e-008             pvth0=3.1474253e-014 k2=0.036557599                lk2=-2.5764511e-013            wk2=-6.8381146e-009 pk2=1.4568607e-019             cit=0.003502                   wcit=-4.54812e-010 voff=-0.084787865               lvoff=-3.4366948e-008            wvoff=-3.5047245e-008 pvoff=2.2627981e-014             eta0=0.1149                     weta0=2.27406e-008 etab=-0.296776                  wetab=-3.9568644e-008            u0=0.014305779 lu0=-1.3779655e-010            wu0=-6.5577506e-010            pu0=1.2484368e-016 ua=1.3962313e-009             lua=-4.9075463e-016            wua=-4.2816443e-016 pua=3.4157648e-022             ub=1.1350954e-018             lub=-2.1750665e-025 wub=-3.1716714e-025            pub=1.7833176e-031             uc=1.4081983e-010 luc=-8.7110118e-022            wuc=-4.9184138e-017            puc=7.717057e-028 vsat=107166.66                  lvsat=4.751519e-008              wvsat=-0.02820266 pvsat=-4.3048762e-014            a0=5.8220252                  la0=-3.0772672e-006 wa0=-3.624027e-006             pa0=3.0676e-012                ags=2.0581851 lags=-9.1922139e-007            wags=-1.4544985e-006            pags=1.7578339e-012 keta=-0.086693153               lketa=5.9823758e-008             wketa=1.0043989e-007 pketa=-9.009458e-014             pclm=0.12974843                 lpclm=1.2028875e-007 wpclm=9.7776966e-008             ppclm=-1.0898179e-013            pdiblc2=0.0010000001 lpdiblc2=-7.522325e-017             wpdiblc2=-1.2629455e-016            ppdiblc2=1.1328622e-022 aigbacc=0.011490979                laigbacc=7.0981367e-011             waigbacc=5.8509496e-010 paigbacc=-8.165897e-017             aigc=0.006029741                laigc=-3.8945985e-011 waigc=-6.362864e-011             paigc=3.3587981e-017             aigsd=0.0048930989 laigsd=6.616015e-012              waigsd=9.284446e-011              paigsd=-5.9941096e-018 tvoff=0.00202911                 ltvoff=-8.92751e-010              wtvoff=-1.1753e-009 ptvoff=1.17201e-015               kt1=-0.23903481                lkt1=2.0586503e-008 wkt1=1.137507e-008              pkt1=-4.8304925e-015            kt2=-0.06 ute=-0.94874906                lute=5.0015989e-013             wute=-2.2763336e-007 pute=-4.5314486e-019            ua1=2.5936535e-009             lua1=-1.1171252e-015 wua1=-1.1014321e-015            pua1=8.383818e-022              ub1=3.1555e-019 lub1=-3.7461953e-026            wub1=-1.2016056e-024            pub1=-8.6348135e-033 uc1=5.2792864e-010             luc1=-3.9378648e-016            wuc1=-5.4529903e-016 puc1=4.8675633e-022             at=90000                      jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)' jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 a0_ff=-0.590147 a0_ss=0.590147                   a0_sf=-0.579086                  a0_fs=0.576346 la0_ff=7.98457e-07                la0_ss=-7.98457e-07               la0_sf=6.98841e-07 la0_fs=-6.74159e-07               wa0_ff=5.04611e-07                wa0_ss=-5.04611e-07 wa0_sf=5.04611e-07                wa0_fs=-5.12149e-07               pa0_ff=-4.52637e-13 pa0_ss=4.52637e-13                pa0_sf=-4.52636e-13               pa0_fs=5.20531e-13 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.2 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.37298288 lvth0=-1.001371e-008             wvth0=-1.1242776e-008            pvth0=3.7804867e-015 k2=0.03801824                 lk2=-1.310453e-009             wk2=-7.3047543e-009 pk2=4.1872144e-016             cit=0.0044953333               wcit=-4.54812e-010 voff=-0.10656722                lvoff=-1.4830864e-008            wvoff=-1.4816225e-008 pvoff=4.4807568e-015             eta0=0.1149                     weta0=2.27406e-008 etab=-0.296776                  wetab=-3.9568644e-008            u0=0.014025923 lu0=1.1323514e-010             wu0=-1.6378346e-009            pu0=1.0057511e-015 ua=1.2499669e-009             lua=-3.5955543e-016            wua=2.3900846e-017 pua=-6.3926071e-023            ub=8.9527423e-019             lub=-2.3870712e-027 wub=-3.4047725e-025            pub=1.9924092e-031             uc=1.358201e-010 luc=4.4838905e-018             wuc=-7.1709276e-017            puc=2.0205821e-023 vsat=107166.72                  lvsat=0                          wvsat=-0.028202708 pvsat=0                          a0=3.5703514                  la0=-1.0575158e-006 wa0=-6.1499941e-007            pa0=3.6850229e-013             ags=0.94853554 lags=7.613426e-008              wags=7.0833905e-007             pags=-1.8223135e-013 keta=-0.0024676667              lketa=-1.5726503e-008            wketa=-3.3883494e-008 pketa=3.0393494e-014             pclm=0.16690838                 lpclm=8.695628e-008 wpclm=1.9087649e-008             ppclm=-3.8397475e-014            pdiblc2=-0.0001229832 lpdiblc2=1.0073159e-009             wpdiblc2=1.1746278e-010             ppdiblc2=-1.0536411e-016 aigbacc=0.011504196                laigbacc=5.9125496e-011             waigbacc=9.6275659e-010 paigbacc=-4.2042145e-016            aigc=0.006013917                laigc=-2.4751794e-011 waigc=-4.9795671e-011            paigc=2.1179808e-017             aigsd=0.004871935 laigsd=2.5600035e-011             waigsd=1.1201896e-010             paigsd=-2.319364e-017 tvoff=0.000591111                ltvoff=3.97131e-010               wtvoff=4.07192e-010 ptvoff=-2.47484e-016              kt1=-0.21856429                lkt1=2.2244429e-009 wkt1=-4.2525255e-009            pkt1=9.1874609e-015             kt2=-0.06 ute=-0.69917216                lute=-2.2386998e-007            wute=-4.5374994e-007 pute=2.0282612e-013             ua1=1.5378978e-009             lua1=-1.701124e-016 wua1=-2.0479568e-016            pua1=3.4098947e-023             ub1=1.3615189e-018 lub1=-9.7569604e-025            wub1=-2.0457691e-024            pub1=7.4857985e-031 uc1=6.0467548e-013             luc1=7.922312e-017              wuc1=-5.2226076e-017 puc1=4.4469886e-023             at=90000                      jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)' jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 lcit=-8.9102e-010 pcit=-8.9026441e-030            u0_ff=9.93332e-05                u0_ss=-4.74399e-06 u0_sf=9.93332e-05                u0_fs=-4.74399e-06               lu0_ff=-8.91019e-11 lu0_ss=4.25488e-12                lu0_sf=-8.91019e-11               lu0_fs=4.25488e-12 wu0_ff=-1.5e-16                   wu0_ss=-6.76991e-11               wu0_sf=-1.5e-16 wu0_fs=-6.76991e-11               pu0_ff=-4.7e-22                   pu0_ss=6.07264e-17 pu0_sf=-4.7e-22                   pu0_fs=6.07264e-17                a0_ff=0.300002 a0_ss=-0.300002                  a0_sf=0.324539                   a0_fs=-0.175225 la0_ff=5.4e-13                    la0_ss=-5.4e-13                   la0_sf=-1.11711e-07 la0_fs=1.5e-13                    wa0_ff=-2.54e-12                  wa0_ss=2.54e-12 wa0_sf=-1.12832e-07               wa0_fs=6.81539e-08                pa0_ff=-5.9e-19 pa0_ss=5.9e-19                    pa0_sf=1.0121e-13                 pa0_fs=-4.7e-19 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.3 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.38899881 lvth0=-2.8545867e-009            wvth0=-2.4024944e-009            pvth0=-1.7111944e-016 k2=0.038912701                lk2=-1.7102772e-009            wk2=-1.2765916e-008 pk2=2.8598607e-015             cit=0.001172894                wcit=5.4183171e-010 voff=-0.13202804                lvoff=-3.4498774e-009            wvoff=-6.3866439e-009 pvoff=7.1273395e-016             eta0=0.1149                     weta0=2.27406e-008 etab=-0.296776                  wetab=-3.9568644e-008            u0=0.012315866 lu0=8.7763024e-010             wu0=1.4134893e-009             pu0=-3.581907e-016 ua=1.3953204e-009             lua=-4.2452844e-016            wua=-1.5964394e-016 pua=1.8118447e-023             ub=4.7549291e-019             lub=1.8525518e-025 wub=2.4840718e-025             pub=-6.3990414e-032            uc=1.4635576e-010 luc=-2.2555224e-019            wuc=-3.7644455e-017            puc=4.9788458e-024 vsat=113315.74                  lvsat=-0.0027486119              wvsat=-0.032128687 pvsat=1.7549127e-009             a0=1.8452868                  la0=-2.864119e-007 wa0=8.9518101e-007             pa0=-3.0654835e-013            ags=3.2956276 lags=-9.7301591e-007            wags=-2.5368272e-006            pags=1.268358e-012 keta=0.019195513                lketa=-2.5409944e-008            wketa=4.4460788e-008 pketa=-4.6264001e-015            pclm=0.26537303                 lpclm=4.2942579e-008 wpclm=-1.043506e-007             ppclm=1.6779424e-014             pdiblc2=0.0013390703 lpdiblc2=3.5377803e-010             wpdiblc2=-2.2588996e-010            ppdiblc2=4.8114561e-017 aigbacc=0.011685459                laigbacc=-2.1899294e-011            waigbacc=-3.035645e-011 paigbacc=2.3500077e-017             aigc=0.0059339944               laigc=1.0973595e-011 waigc=2.0396692e-011             paigc=-1.0196179e-017            aigsd=0.0049444082 laigsd=-6.795514e-012             waigsd=3.4419503e-011             paigsd=1.149332e-017 tvoff=0.00197337                 ltvoff=-2.20739e-010              wtvoff=-5.56614e-010 ptvoff=1.83337e-016               kt1=-0.20541505                lkt1=-3.6532665e-009 wkt1=2.4341346e-008             pkt1=-3.5939995e-015            kt2=-0.055448718 ute=-1.3376775                 lute=6.1541909e-008             wute=2.0720495e-007 pute=-9.2620716e-014            ua1=1.3809769e-009             lua1=-9.9968751e-017 wua1=-3.2000945e-016            pua1=8.5599506e-023             ub1=-1.4228015e-018 lub1=2.6889515e-025             wub1=-2.1969562e-025            pub1=-6.7675009e-032 uc1=7.9091999e-011             luc1=4.4139287e-017             wuc1=1.5898934e-016 puc1=-4.9943405e-023            at=71035.665 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=5.9411038e-010             pcit=-4.4549974e-016            lkt2=-2.0344231e-009 lat=0.0084770576               wat=0.050094971                pat=-2.2392452e-008 u0_ff=3.65388e-05                u0_ss=-4.0738e-05                u0_sf=-8.97423e-06 u0_fs=-4.0738e-05                lu0_ff=-6.1033e-11                lu0_ss=2.03444e-11 lu0_sf=-4.06886e-11               lu0_fs=2.03444e-11                wu0_ff=6e-17 wu0_ss=6.81541e-11                wu0_sf=6e-17                      wu0_fs=6.81541e-11 pu0_ff=-1.17e-22                  pu0_ss=-7e-24                     pu0_sf=1.83e-22 pu0_fs=-7e-24                     a0_ff=0.299997                   a0_ss=-0.299997 a0_sf=-0.039497                  a0_fs=-0.015453                  la0_ff=-4e-14 la0_ss=4e-14                      la0_sf=5.10123e-08                la0_fs=-7.14177e-08 wa0_ff=-2.7e-12                   wa0_ss=2.7e-12                    wa0_sf=2.16985e-07 wa0_fs=-7.65994e-08               pa0_ff=1.5e-19                    pa0_ss=-1.5e-19 pa0_sf=-4.62182e-14               pa0_fs=6.47046e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.4 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.39832837 lvth0=-8.6739128e-010            wvth0=-2.6534294e-009            pvth0=-1.1767028e-016 k2=0.037031841                lk2=-1.309654e-009             wk2=4.7834789e-009 pk2=-8.7816039e-016            cit=0.0047985641               wcit=-1.6571428e-009 voff=-0.13067548                lvoff=-3.7379743e-009            wvoff=-6.1804621e-009 pvoff=6.6881723e-016             eta0=0.1149                     weta0=2.27406e-008 etab=-0.29678516                wetab=-3.9558921e-008            u0=0.016299128 lu0=2.9195618e-011             wu0=-6.4081056e-010            pu0=7.9375176e-017 ua=-2.1523823e-010            lua=-8.1479455e-017            wua=-2.3353304e-016 pua=3.3856825e-023             ub=1.4186773e-018             lub=-1.5643099e-026 wub=9.439888e-026              pub=-3.1186647e-032            uc=2.1326912e-010 luc=-1.4478098e-017            wuc=-2.3177477e-017            puc=1.8973794e-024 vsat=94150.336                  lvsat=0.0013336184               wvsat=-0.018684898 pvsat=-1.1086145e-009            a0=0.28768123                 la0=4.5358083e-008 wa0=2.1312947e-006             pa0=-5.6984057e-013            ags=-3.5321208 lags=4.8129451e-007             wags=5.7778871e-006             pags=-5.0267618e-013 keta=-0.068160084               lketa=-6.8032021e-009            wketa=-6.1969637e-009 pketa=6.1637011e-015             pclm=0.49208413                 lpclm=-5.346884e-009 wpclm=-2.4073623e-008            ppclm=-3.1957295e-016            pdiblc2=0.0023095238 lpdiblc2=1.4707143e-010             wpdiblc2=0                          ppdiblc2=0 aigbacc=0.011312385                laigbacc=5.7565583e-011             waigbacc=7.8574087e-010 paigbacc=-1.5032865e-016            aigc=0.0059853203               laigc=4.1184397e-014 waigc=-5.7672647e-012            paigc=-4.6232559e-018            aigsd=0.0048068453 laigsd=2.2505387e-011             waigsd=9.8668277e-011             paigsd=-2.1916694e-018 tvoff=0.000818232                ltvoff=2.53055e-011               wtvoff=4.71945e-010 ptvoff=-3.57461e-017              kt1=-0.2051248                 lkt1=-3.7150907e-009 wkt1=-1.9214952e-008            pkt1=5.6834918e-015             kt2=-0.065 ute=-0.87526506                lute=-3.6951939e-008            wute=-3.8481001e-007 pute=3.347847e-014              ua1=1.4463704e-009             lua1=-1.1389757e-016 wua1=-6.7191948e-017            pua1=3.1749377e-023             ub1=-2.2166158e-019 lub1=1.3052359e-026             wub1=-7.6965998e-025            pub1=4.94674e-032 uc1=3.6475417e-010             luc1=-1.6706755e-017            wuc1=-1.1229924e-016 puc1=7.8410624e-024             at=131066.7                   jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)' jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 lcit=-1.7815736e-010 pcit=2.2881834e-017             lat=-0.0043095521              wat=-0.063364713 pat=1.7744607e-009             letab=1.9511849e-012             petab=-2.0709098e-018 u0_ff=-0.000388097               u0_ss=-4.54983e-05               u0_sf=-0.000338096 u0_fs=9.25967e-05                lu0_ff=2.94142e-11                lu0_ss=2.13584e-11 lu0_sf=2.94143e-11                lu0_fs=-8.05592e-12               wu0_ff=-6e-17 wu0_ss=1.15213e-10                wu0_sf=-2.5e-16                   wu0_fs=1.15212e-10 pu0_ff=1.8e-23                    pu0_ss=-1.00235e-17               pu0_sf=-5e-24 pu0_fs=-1.00235e-17               vsat_ff=2421.84                    vsat_ss=-2421.84 lvsat_ff=-0.000515852               lvsat_ss=0.000515852                wvsat_ff=-0.00156862 wvsat_ss=0.00156862                 pvsat_ff=3.34115e-10                pvsat_ss=-3.34115e-10 a0_ff=0.0918189                  a0_ss=-0.0918189                 a0_sf=0.0959121 a0_fs=-0.592933                  la0_ff=4.43416e-08                la0_ss=-4.43416e-08 la0_sf=2.21708e-08                la0_fs=5.15852e-08                wa0_ff=3.13722e-07 wa0_ss=-3.13722e-07               wa0_sf=1.56862e-07                wa0_fs=3.84039e-07 pa0_ff=-6.68236e-14               pa0_ss=6.68236e-14                pa0_sf=-3.34115e-14 pa0_fs=-3.34115e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.5 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.38194061 lvth0=-2.2931268e-009            wvth0=-1.9193531e-008            pvth0=1.3213186e-015 k2=0.056519861                lk2=-3.0051118e-009            wk2=-7.3352766e-009 pk2=1.7617133e-016             cit=4.7046082e-005             wcit=-1.2159155e-009 voff=-0.13064829                lvoff=-3.7403391e-009            wvoff=-5.2946143e-009 pvoff=5.9174848e-016             eta0=0.143375                   weta0=-9.47525e-009 etab=-0.51824888                wetab=-1.4480352e-007            u0=0.017195353 lu0=-4.8775948e-011            wu0=3.6205499e-010             pu0=-7.8741272e-018 ua=-1.655312e-009             lua=4.3806961e-017             wua=6.1182572e-016 pua=-3.9689387e-023            ub=2.1428133e-018             lub=-7.8642932e-026 wub=-8.8342507e-025            pub=5.3884037e-032             uc=2.3275161e-010 luc=-1.6173074e-017            wuc=-8.724216e-017             puc=7.4710069e-024 vsat=119304.62                  lvsat=-0.0008548044              wvsat=-0.062892065 pvsat=2.7374091e-009             a0=18.007918                  la0=-1.4963025e-006 wa0=-1.6094578e-005            pa0=1.0158103e-012             ags=2 lags=0                          wags=0                          pags=0 keta=-0.024789165               lketa=-1.0576472e-008            wketa=-4.6670641e-008 pketa=9.684911e-015              pclm=0.66556525                 lpclm=-2.0439742e-008 wpclm=-1.6943212e-007            ppclm=1.2326616e-014             pdiblc2=0.0025833333 lpdiblc2=1.2325e-010                wpdiblc2=0                          ppdiblc2=0 aigbacc=0.011765724                laigbacc=1.8125036e-011             waigbacc=-1.1726411e-009 paigbacc=2.0050576e-017             aigc=0.0061689783               laigc=-1.5937064e-011 waigc=-1.336876e-010             paigc=6.5058133e-018             aigsd=0.004914434 laigsd=1.3145172e-011             waigsd=1.5570409e-010             paigsd=-7.153785e-018 tvoff=0.00165215                 ltvoff=-4.72449e-011              wtvoff=-7.44821e-010 ptvoff=7.01125e-017               kt1=-0.25751409                lkt1=8.4277761e-010 wkt1=7.3577103e-008             pkt1=-2.389417e-015             kt2=-0.036489374 ute=-1.4416667                 lute=1.2325e-008                ua1=5.952099e-011 lua1=6.7583255e-018             wua1=6.2608814e-016             pua1=-2.8565991e-023 ub1=-5.0315439e-019            lub1=3.7542234e-026             wub1=-4.1174738e-025 pub1=1.8329004e-032             uc1=9.1324375e-011             luc1=7.0816369e-018 wuc1=4.4059913e-018             puc1=-2.3122926e-024            at=97455.356 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=2.3522471e-010             pcit=-1.5504942e-017            lkt2=-2.4804245e-009 lat=-0.0013853654              wat=-0.076715293               pat=2.9359612e-009 letab=1.9269294e-008             petab=9.1542096e-015             leta0=-2.477325e-009 peta0=2.802779e-015              wkt2=-3.2248127e-008            pkt2=2.805587e-015 u0_ff=-0.000120833               u0_ss=0.000483331                lu0_ff=6.16251e-12 lu0_ss=-2.465e-11                 wu0_ff=-2e-16                     wu0_ss=-1.2e-15 pu0_ff=-3.3e-23                   pu0_ss=3.2e-23                    vsat_ff=-3507.47 vsat_ss=3507.47                    lvsat_ff=-1.6e-10                   lvsat_ss=1.6e-10 wvsat_ff=0.0022718                  wvsat_ss=-0.0022718                 pvsat_ff=-3.4e-16 pvsat_ss=3.4e-16                    a0_ff=1.45362                    a0_ss=-1.45362 a0_sf=0.847641                   la0_ff=-7.41346e-08               la0_ss=7.41346e-08 la0_sf=-4.32298e-08               wa0_ff=-1.09803e-06               wa0_ss=1.09803e-06 wa0_sf=-5.49016e-07               pa0_ff=5.59995e-14                pa0_ss=-5.59995e-14 pa0_sf=2.79998e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.6 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.4254328 lvth0=-7.502483e-011             wvth0=3.7721233e-008             pvth0=-1.5813344e-015 k2=0.070438433                lk2=-3.7149589e-009            wk2=-3.5599972e-008 pk2=1.6176708e-015             cit=0.0034248233               wcit=-8.793924e-009 voff=-0.16832318                lvoff=-1.8189199e-009            wvoff=5.1879603e-008 pvoff=-2.3241366e-015            eta0=-0.1806192                 weta0=3.1970252e-007 etab=-0.65353655                wetab=2.1131378e-007             u0=0.016717525 lu0=-2.4406769e-011            wu0=-3.4730885e-010            pu0=2.8303428e-017 ua=-1.6072314e-009            lua=4.1354853e-017             wua=-2.1273533e-017 pua=-7.4013251e-024            ub=2.1199616e-018             lub=-7.7477491e-026 wub=-6.5916263e-025            pub=4.2446652e-032             uc=3.2223598e-010 luc=-2.0736777e-017            wuc=-2.7175714e-016            puc=1.6881271e-023 vsat=72386.501                  lvsat=0.0015380197               wvsat=-0.017067937 pvsat=4.0037858e-010             a0=-23.174685                 la0=6.0401024e-007 wa0=2.6766335e-005             pa0=-1.1700962e-012            ags=2 lags=0                          wags=0                          pags=0 keta=-0.46795513                lketa=1.2024992e-008             wketa=2.8270205e-007 pketa=-7.1130962e-015            pclm=0.40399267                 lpclm=-7.09954e-009 wpclm=-5.7617669e-008            ppclm=6.6240793e-015             pdiblc2=0.00033333333 lpdiblc2=2.38e-010                  wpdiblc2=0                          ppdiblc2=0 aigbacc=0.014339033                laigbacc=-1.1311371e-010            waigbacc=-4.0285482e-009 paigbacc=1.6570184e-016             aigc=0.0061846241               laigc=-1.6735002e-011 waigc=-1.5961876e-010            paigc=7.8283023e-018             aigsd=0.0050901352 laigsd=4.1844132e-012             waigsd=5.3816289e-011             paigsd=-1.9575072e-018 tvoff=-0.00245762                ltvoff=1.62353e-010               wtvoff=3.53827e-009 ptvoff=-1.48325e-016              kt1=-0.21936481                lkt1=-1.1028352e-009 wkt1=4.8679211e-009             pkt1=1.1147513e-015             kt2=-0.20237588 ute=-1.2                       ua1=1.0400629e-009             lua1=-4.3249312e-017 wua1=-2.5407651e-016            pua1=1.6322406e-023             ub1=-1.7141262e-018 lub1=9.9301794e-026             wub1=1.2811524e-024             pub1=-6.8008884e-032 uc1=4.8302e-010                luc1=-1.289484e-017             wuc1=-2.3195412e-016 puc1=9.742073e-024              at=92413.924 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=6.2958071e-011             pcit=3.7097349e-016             lkt2=5.9797873e-009 lat=-0.0011282524              wat=-0.04591329                pat=1.3650591e-009 letab=2.6168966e-008             petab=-9.0077728e-015            leta0=1.4046379e-008 peta0=-1.3985287e-014            wkt2=1.2899255e-007             pkt2=-5.4176875e-015 vsat_ff=-3507.49                   vsat_ss=3507.49                    lvsat_ff=-3.97e-09 lvsat_ss=3.97e-09                   wvsat_ff=0.00227181                 wvsat_ss=-0.00227181 pvsat_ff=-5.2e-16                   pvsat_ss=5.2e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.7 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=9e-007                     wmax=1.3501e-06                 vth0=-0.38934128 lvth0=-1.5908686e-009            wvth0=6.1807116e-009             pvth0=-2.566325e-016 k2=-0.0055783145              lk2=-5.2225555e-010            wk2=7.6048081e-009 pk2=-1.9692997e-016            cit=-0.015251522               wcit=2.758255e-009 voff=-0.13530613                lvoff=-3.2056361e-009            wvoff=1.064163e-008 pvoff=-5.9214173e-016            eta0=0.21383587                 weta0=-1.0366682e-007 etab=-0.14646132                wetab=-2.9521035e-008            u0=0.014756431 lu0=5.7959185e-011             wu0=8.1849226e-010             pu0=-2.0660218e-017 ua=-1.5792903e-010            lua=-1.9515848e-017            wua=-1.2128607e-015 pua=4.2645335e-023             ub=-8.0674532e-019            lub=4.5444198e-026 wub=2.1854156e-024             pub=-7.7025633e-032            uc=-6.0842762e-010 luc=1.8351094e-017             wuc=6.0008644e-016             puc=-1.973616e-023 vsat=106966.41                  lvsat=8.5663606e-005             wvsat=-0.01904671 pvsat=4.8348705e-010             a0=-4.7321433                 la0=-1.7057651e-007 wa0=2.8447325e-005             pa0=-1.2406978e-012            ags=2 lags=0                          wags=0                          pags=0 keta=-0.5774873                 lketa=1.6625343e-008             wketa=6.3294729e-007 pketa=-2.1823396e-014            pclm=0.0086744479               lpclm=9.5038252e-009 wpclm=5.0389807e-007             ppclm=-1.6959582e-014            pdiblc2=0.00787 lpdiblc2=-7.854e-011                wpdiblc2=-8.33822e-009              ppdiblc2=3.5020524e-016 aigbacc=0.0077471602               laigbacc=1.6374495e-010             waigbacc=5.7916309e-009 paigbacc=-2.4674568e-016            aigc=0.0061666962               laigc=-1.598203e-011 waigc=-1.9817719e-010            paigc=9.4477564e-018             aigsd=0.0050206882 laigsd=7.1011848e-012             waigsd=1.603945e-010              paigsd=-6.4337921e-018 tvoff=0.00419159                 ltvoff=-1.16914e-010              wtvoff=-2.03238e-009 ptvoff=8.56423e-017               kt1=-0.14186569                lkt1=-4.3577984e-009 wkt1=-3.8600102e-008            pkt1=2.9404083e-015             kt2=-0.14272943 ute=-1.2                       ua1=4.8599504e-009             lua1=-2.0368459e-016 wua1=-2.3635085e-015            pua1=1.0491855e-022             ub1=-7.8750479e-018 lub1=3.5806051e-025             wub1=4.6940948e-024             pub1=-2.1135246e-031 uc1=3.41e-010                  luc1=-6.93e-018                 at=66005.353 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=8.4736458e-010             pcit=-1.1421803e-016            lkt2=3.4746363e-009 lat=-1.9092421e-005            wat=-0.023998346               pat=4.4463139e-010 letab=4.8718064e-009             petab=1.1072893e-015             leta0=-2.5207336e-009 peta0=3.7962248e-015             wkt2=4.1732857e-008             pkt2=-1.7527804e-015 vth0_ss=-0.0110549                 vth0_mc=0.0200298                  lvth0_ss=4.64306e-10 lvth0_mc=-8.41235e-10               wvth0_ss=1.66597e-08                wvth0_mc=4.16497e-08 pvth0_ss=-6.99709e-16               pvth0_mc=-1.74927e-15               cit_mc=0.0110549 wcit_mc=-1.66597e-08               voff_mc=0.0293334                  lvoff_mc=-1.232e-09 wvoff_mc=-1.2e-14                   pvoff_mc=2.5e-21                    u0_mc=0.00221098 lu0_mc=-9.28612e-11               wu0_mc=-3.33195e-09               pu0_mc=1.39942e-16 vsat_ff=-10840.9                   vsat_sf=4421.96                    vsat_ss=16368.3 vsat_mc=22109.8                    lvsat_ff=0.000308                   lvsat_sf=-0.000185722 lvsat_ss=-0.000540153               lvsat_mc=-0.000928612               wvsat_ff=0.00227174 wvsat_sf=-0.0066639                 wvsat_ss=-0.0106016                 wvsat_mc=-0.0333195 pvsat_ff=6.9e-16                    pvsat_sf=2.79884e-10                pvsat_ss=3.49854e-10 pvsat_mc=1.39942e-09                lcit_mc=-4.64306e-10               pcit_mc=6.99709e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model pch_lvt_mac.8 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.40801819 lvth0=1.7841372e-008             wvth0=1.3025935e-008             pvth0=-1.4752688e-014 k2=0.036904273                lk2=-2.0594565e-013            wk2=-7.1522015e-009 pk2=9.884636e-020              cit=0.0028483333               wcit=1.3741e-010 voff=-0.13393821                lvoff=-1.9794243e-009            wvoff=9.4829678e-009 pvoff=-6.7151152e-015            eta0=0.14                       weta0=0 etab=-0.38452433                wetab=3.9931346e-008             u0=0.012533925 lu0=0                          wu0=9.4952509e-010             pu0=0 ua=7.9941658e-010             lua=3.393733e-017              wua=1.1254972e-016 pua=-1.3379443e-022            ub=8.0013337e-019             lub=-1.1970515e-026 wub=-1.3691543e-026            pub=-7.8839843e-033            uc=1.2355241e-010 luc=-3.5044404e-023            wuc=-3.3539859e-017            puc=1.4238257e-029 vsat=71546.595                  lvsat=0                          wvsat=0.0040691223 pvsat=0                          a0=0.3119247                  la0=1.9129571e-006 wa0=1.3681241e-006             pa0=-1.4535432e-012            ags=-0.1453673 lags=2.0796338e-006             wags=5.4191995e-007             pags=-9.5912885e-013 keta=0.015321922                lketa=-9.9706264e-008            wketa=8.0142308e-009 pketa=5.443962e-014              pclm=0.21896956                 lpclm=-5.0148834e-013 wpclm=1.6942623e-008             ppclm=2.7381263e-019             pdiblc2=0.00094650562 lpdiblc2=4.8128778e-010             wpdiblc2=4.8465856e-011             ppdiblc2=-4.3604668e-016 aigbacc=0.011817137                laigbacc=-3.9936587e-011            waigbacc=2.8959578e-010 paigbacc=1.8832696e-017             aigc=0.0059328547               laigc=3.2683628e-011 waigc=2.4150422e-011             paigc=-3.1308448e-017            aigsd=0.0049646534 laigsd=-1.511107e-017             waigsd=2.8016015e-011             paigsd=1.3690636e-023 tvoff=0.00120583                 ltvoff=3.7261e-010                wtvoff=-4.29417e-010 ptvoff=2.55939e-017               kt1=-0.20858041                lkt1=-1.2063147e-009 wkt1=-1.6216616e-008            pkt1=1.4913801e-014             kt2=-0.044833333 ute=-1.4080867                 wute=1.8852652e-007             ua1=5.1059056e-010 lua1=1.3341372e-016             wua1=7.8582291e-016             pua1=-2.9460651e-022 ub1=-1.6441606e-018            lub1=1.512629e-025              wub1=5.7389215e-025 pub1=-1.7961953e-031            uc1=-7.2296372e-010            luc1=4.5627136e-016 wuc1=5.8800945e-016             puc1=-2.8339607e-022            at=105166.67 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' wat=-0.013741                  wkt2=-1.3741e-008               a0_ff=0.13526 a0_ss=-0.13526                   a0_sf=0.146321                   a0_fs=-0.157381 la0_ff=1.47772e-07                la0_ss=-1.47772e-07               la0_sf=4.81507e-08 la0_fs=5.14712e-08                wa0_ff=-1.52608e-07               wa0_ss=1.52608e-07 wa0_sf=-1.52608e-07               wa0_fs=1.52608e-07                pa0_ff=1.36889e-13 pa0_ss=-1.36889e-13               pa0_sf=1.36889e-13                pa0_fs=-1.3689e-13 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.9 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.38189812 lvth0=-5.588325e-009             wvth0=-3.1655656e-009            pvth0=-2.2891193e-016 k2=0.03763138                 lk2=-6.5242147e-010            wk2=-6.9542594e-009 pk2=-1.7745517e-016            cit=0.0035686788               wcit=3.8473701e-010 voff=-0.12531713                lvoff=-9.712529e-009             wvoff=2.1711949e-009 pvoff=-1.5645486e-016            eta0=0.14                       weta0=0 etab=-0.38452433                wetab=3.9931346e-008             u0=0.010222147 lu0=2.0736648e-009             wu0=1.8083859e-009             pu0=-7.7039812e-016 ua=1.2728525e-009             lua=-3.9073467e-016            wua=3.1664936e-018 pua=-3.5677678e-023            ub=4.7043422e-019             lub=2.8376962e-025 wub=4.4427804e-026             pub=-6.0017039e-032            uc=8.0419755e-011 luc=3.868996e-017              wuc=-2.1516567e-017            puc=-1.0784879e-023 vsat=71546.595                  lvsat=0                          wvsat=0.0040691223 pvsat=0                          a0=3.1156986                  la0=-6.0202814e-007 wa0=-2.03084e-007              pa0=-4.4169512e-014            ags=2.133797 lags=3.5223449e-008             wags=-3.6550781e-007            pags=-1.4516615e-013 keta=-0.13076556                lketa=3.1334203e-008             wketa=8.2354393e-008 pketa=-1.2243506e-014            pclm=0.085573542                lpclm=1.1965572e-007 wpclm=9.2777008e-008             ppclm=-6.802317e-014             pdiblc2=0.00096956294 lpdiblc2=4.6060536e-010             wpdiblc2=-8.7238403e-010            ppdiblc2=3.8995566e-016 aigbacc=0.011913006                laigbacc=-1.2593188e-010            waigbacc=5.9237411e-010 paigbacc=-2.5275946e-016            aigc=0.005979511                laigc=-9.1670686e-012 waigc=-1.862382e-011             paigc=7.0600462e-018             aigsd=0.0049646534 laigsd=-8.9101959e-018            waigsd=2.801603e-011              paigsd=2.6004101e-030 tvoff=0.00184914                 ltvoff=-2.04434e-010              wtvoff=-7.32582e-010 ptvoff=2.97534e-016               kt1=-0.21753013                lkt1=6.821581e-009 wkt1=-5.1894734e-009            pkt1=5.0224538e-015             kt2=-0.044833333 ute=-1.4748268                 lute=5.9865925e-008             wute=2.489932e-007 pute=-5.4238608e-014            ua1=3.8464628e-010             lua1=2.4638574e-016 wua1=8.4005017e-016             pua1=-3.4324836e-022            ub1=-1.3095745e-018 lub1=-1.4886077e-025            wub1=3.7424151e-025             pub1=-5.3290594e-034 uc1=-3.9376282e-010            luc1=1.6097815e-016             wuc1=3.0507087e-016 puc1=-2.9600169e-023            at=120232.22 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=-6.4614988e-010            pcit=-2.2185233e-016            lat=-0.013513803 wat=-0.027390393               pat=1.2243506e-008             wkt2=-1.3741e-008 u0_ff=2.40057e-05                u0_ss=-4.93354e-05               u0_sf=9.93334e-05 u0_fs=-4.93354e-05               lu0_ff=-2.15329e-11               lu0_ss=4.4254e-11 lu0_sf=-8.9102e-11                lu0_fs=4.4254e-11                 wu0_ff=6.82469e-11 wu0_ss=-2.72989e-11               wu0_sf=-7e-17                     wu0_fs=-2.72989e-11 pu0_ff=-6.12176e-17               pu0_ss=2.44871e-17                pu0_sf=-6e-23 pu0_fs=2.44871e-17                a0_ff=0.300003                   a0_ss=-0.300003 a0_sf=0.199999                   a0_fs=-0.130131                  la0_ff=-1e-13 la0_ss=1e-13                      la0_sf=-7e-14                     la0_fs=2.70276e-08 wa0_ff=2e-13                      wa0_ss=-2e-13                     wa0_sf=1.3e-13 wa0_fs=2.72987e-08                pa0_ff=1.7e-19                    pa0_ss=-1.7e-19 pa0_sf=1.2e-19                    pa0_fs=-2.44871e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.10 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.37971545 lvth0=-6.5639819e-009            wvth0=-1.0813227e-008            pvth0=3.1895926e-015 k2=0.031437453                lk2=2.1162639e-009             wk2=-5.9933412e-009 pk2=-6.0698562e-016            cit=0.0029211239               wcit=-1.0420645e-009 voff=-0.13727429                lvoff=-4.36768e-009              wvoff=-1.6335433e-009 pvoff=1.5442631e-015             eta0=0.14                       weta0=0 etab=-0.38452433                wetab=3.9931346e-008             u0=0.013996277 lu0=3.8662879e-010             wu0=-1.0896252e-010            pu0=8.6656609e-017 ua=1.4424706e-009             lua=-4.6655397e-016            wua=-2.0236204e-016 pua=5.6193576e-023             ub=8.0193967e-019             lub=1.3558668e-025 wub=-4.7353589e-026            pub=-1.8990756e-032            uc=1.6786857e-010 luc=-3.9966107e-019            wuc=-5.7135061e-017            puc=5.1365884e-024 vsat=75444.304                  lvsat=-0.001742276               wvsat=0.0021828307 pvsat=8.4317234e-010             a0=3.3188053                  la0=-6.9281683e-007 wa0=-4.398268e-007             pa0=6.1654519e-014             ags=1.9509859 lags=1.1694e-007                wags=-1.3185818e-006            pags=2.8085793e-013 keta=0.028310897                lketa=-3.9772971e-008            wketa=3.620225e-008 pketa=8.3865022e-015             pclm=0.24726168                 lpclm=4.7381124e-008 wpclm=-8.7941722e-008            ppclm=1.2758102e-014             pdiblc2=0.0010897436 lpdiblc2=4.0688462e-010             wpdiblc2=0                          ppdiblc2=0 aigbacc=0.011585506                laigbacc=2.0460851e-011             waigbacc=6.0201291e-011 paigbacc=-1.4878214e-017            aigc=0.0059730765               laigc=-6.2908786e-012 waigc=-1.5011712e-011            paigc=5.4454342e-018             aigsd=0.0049836165 laigsd=-8.4765188e-012            waigsd=-1.1032314e-012            paigsd=1.301631e-017 tvoff=0.0013998                  ltvoff=-3.58144e-012              wtvoff=-3.69642e-011 ptvoff=-1.34076e-017              kt1=-0.18985611                lkt1=-5.5487046e-009 wkt1=1.0244948e-008             pkt1=-1.8767326e-015            kt2=-0.033379273 ute=-1.2400711                 lute=-4.5069869e-008            wute=1.1877359e-007 pute=3.9695551e-015             ua1=8.1074905e-010             lua1=5.5917799e-017 wua1=1.9661694e-016             pua1=-5.5633708e-023            ub1=-2.1017933e-018 lub1=2.05261e-025               wub1=3.9547095e-025             pub1=-1.0022464e-032 uc1=-1.4962919e-010            luc1=5.1850419e-017             wuc1=3.6621074e-016 puc1=-5.6929691e-023            at=122744.75 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=-3.5669283e-010            pcit=4.1592796e-016             lkt2=-5.1199647e-009 lat=-0.014636904               wat=0.0032465382               pat=-1.4512026e-009 wkt2=-1.9994917e-008            pkt2=2.7955007e-015             u0_ff=0.000181399 u0_ss=4.15378e-06                u0_sf=-8.97478e-06               u0_fs=4.15378e-06 lu0_ff=-9.18882e-11               lu0_ss=2.03441e-11                lu0_sf=-4.06891e-11 lu0_fs=2.03441e-11                wu0_ff=-1.31245e-10               wu0_ss=2.74823e-11 wu0_sf=-3.3e-16                   wu0_fs=2.74823e-11                pu0_ff=2.7955e-17 pu0_ss=-1.5e-23                   pu0_sf=1.5e-23                    pu0_fs=-1.5e-23 a0_ff=0.369023                   a0_ss=-0.299996                  a0_sf=0.200001 a0_fs=-0.0420559                 la0_ff=-3.08559e-08               la0_ss=5e-13 la0_sf=-6.7e-13                   la0_fs=-1.23425e-08               wa0_ff=-6.25392e-08 wa0_ss=0.0                        wa0_sf=3.3e-13                    wa0_fs=-5.24977e-08 pa0_ff=2.7955e-14                 pa0_ss=-5e-20                     pa0_sf=3e-20 pa0_fs=1.1182e-14 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.11 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.40499676 lvth0=-1.1790612e-009            wvth0=3.3881345e-009             pvth0=1.6470263e-016 k2=0.055736417                lk2=-3.0594152e-009            wk2=-1.2162866e-008 pk2=7.0712324e-016             cit=0.0013356844               wcit=1.4802262e-009 voff=-0.14327972                lvoff=-3.0885237e-009            wvoff=5.2389832e-009 pvoff=8.0414981e-017             eta0=0.14                       weta0=0 etab=-0.38451985                wetab=3.9928704e-008             u0=0.015111015 lu0=1.4918957e-010             wu0=4.3561944e-010             pu0=-2.9339348e-017 ua=-6.0739853e-010            lua=-2.9931844e-017            wua=1.2176419e-016 pua=-1.2845311e-023            ub=1.7355527e-018             lub=-6.3272887e-026 wub=-1.9269019e-025            pub=1.1965941e-032             uc=2.2613526e-010 luc=-1.2810465e-017            wuc=-3.4834198e-017            puc=3.8650441e-025 vsat=68587.447                  lvsat=-0.00028176534             wvsat=0.00447508 pvsat=3.5492325e-010             a0=3.6185527                  la0=-7.5666301e-007 wa0=-8.8647481e-007            pa0=1.5679054e-013             ags=2.8452381 lags=-7.3535714e-008            wags=0                          pags=0 keta=-0.18983333                lketa=6.69175e-009               wketa=1.04039e-007 pketa=-6.0627255e-015            pclm=0.52106998                 lpclm=-1.0940044e-008 wpclm=-5.0334809e-008            ppclm=4.7478299e-015             pdiblc2=0.0023095238 lpdiblc2=1.4707143e-010             wpdiblc2=0                          ppdiblc2=0 aigbacc=0.012079436                laigbacc=-8.4746167e-011            waigbacc=9.0792804e-011 paigbacc=-2.1394206e-017            aigc=0.0059718766               laigc=-6.0352852e-012 waigc=6.4127415e-012             paigc=8.8202551e-019             aigsd=0.0048119264 laigsd=2.8093478e-011             waigsd=9.4064794e-011             paigsd=-7.2544795e-018 tvoff=0.00139082                 ltvoff=-1.66874e-012              wtvoff=-4.68242e-011 ptvoff=-1.13074e-017              kt1=-0.2399163                 lkt1=5.114115e-009 wkt1=1.230615e-008              pkt1=-2.3157685e-015            kt2=-0.055343167 ute=-1.4516668                 lute=1.4707143e-014             wute=1.3741e-007 pute=-4.715599e-028             ua1=1.5420831e-009             lua1=-9.9856344e-017 wua1=-1.5390763e-016            pua1=1.9028025e-023             ub1=-1.6531028e-018 lub1=1.0968993e-025             wub1=5.2722577e-025             pub1=-3.808624e-032 uc1=9.4688988e-011             luc1=-1.8935446e-019            wuc1=1.3237981e-016 puc1=-7.1237025e-024            at=69493.237 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=-1.8994224e-011            pcit=-1.2131997e-016            lkt2=-4.416555e-010 lat=-0.0032943313              wat=-0.0075791579              pat=8.5467068e-010 letab=-9.5580496e-013            petab=5.6282302e-019             wkt2=-8.749091e-009 pkt2=4.0013988e-016             u0_ff=-0.000335734               u0_ss=3.03877e-05 u0_sf=-0.000338095               u0_fs=0.000168484                lu0_ff=1.82613e-11 lu0_ss=1.47562e-11                lu0_sf=2.94143e-11                lu0_fs=-1.46582e-11 wu0_ff=-4.74388e-11               wu0_ss=4.64575e-11                wu0_sf=3.3e-16 wu0_fs=4.64575e-11                pu0_ff=1.01045e-17                pu0_ss=-4.04183e-18 pu0_sf=-3e-23                     pu0_fs=-4.04183e-18               vsat_ff=690.478 vsat_ss=-690.478                   lvsat_ff=-0.000147072               lvsat_ss=0.000147072 wvsat_ff=3.3e-10                    wvsat_ss=-3.3e-10                   pvsat_ff=1.5e-16 pvsat_ss=-1.5e-16                   a0_ff=0.309901                   a0_ss=-0.438095 a0_sf=0.269047                   a0_fs=-0.169048                  la0_ff=-1.82614e-08 la0_ss=2.94143e-08                la0_sf=-1.47072e-08               la0_fs=1.47072e-08 wa0_ff=1.16144e-07                wa0_ss=3.33e-13                   wa0_sf=-6.33e-13 wa0_fs=-3.3e-13                   pa0_ff=-1.01045e-14               pa0_ss=1.5e-20 pa0_sf=-1.5e-20                   pa0_fs=-1.5e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.12 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.41504109 lvth0=-3.0520465e-010            wvth0=1.0795508e-008             pvth0=-4.7973889e-016 k2=0.060015407                lk2=-3.4316874e-009            wk2=-1.0502241e-008 pk2=5.6264881e-016             cit=-0.0015528093              wcit=2.3355349e-010 voff=-0.14681436                lvoff=-2.7810096e-009            wvoff=9.3518457e-009 pvoff=-2.7740405e-016            eta0=0.13291667                 weta0=0 etab=-0.75738294                wetab=7.1851938e-008             u0=0.019074904 lu0=-1.9566882e-010            wu0=-1.3408192e-009            pu0=1.2521081e-016 ua=-7.2420192e-010            lua=-1.9769949e-017            wua=-2.3175999e-016 pua=1.7911293e-023             ub=1.0984255e-018             lub=-7.8428235e-027 wub=6.279029e-026              pub=-1.0260861e-032            uc=2.389245e-010 luc=-1.3923129e-017            wuc=-9.2834797e-017            puc=5.4325565e-024 vsat=32129.026                  lvsat=0.0028901173               wvsat=0.016089025 pvsat=-6.5548993e-010            a0=-1.5213642                 la0=-3.0949025e-007 wa0=1.5989517e-006             pa0=-5.9441565e-014            ags=2 lags=0                          wags=0                          pags=0 keta=-0.14268272                lketa=2.5896469e-009             wketa=6.0140922e-008 pketa=-2.2435927e-015            pclm=0.54094283                 lpclm=-1.2668982e-008 wpclm=-5.6524207e-008            ppclm=5.2863075e-015             pdiblc2=0.0025833333 lpdiblc2=1.2325e-010                wpdiblc2=0                          ppdiblc2=0 aigbacc=0.010346455                laigbacc=6.6023166e-011             waigbacc=1.1321721e-010 paigbacc=-2.3345129e-017            aigc=0.0059922017               laigc=-7.8035717e-012 waigc=2.6472006e-011             paigc=-8.6313046e-019            aigsd=0.0050779623 laigsd=4.9483537e-012             waigsd=7.5474172e-012             paigsd=2.7253231e-019 tvoff=0.00190504                 ltvoff=-4.64056e-011              wtvoff=-9.73945e-010 ptvoff=6.93521e-017               kt1=-0.11108963                lkt1=-6.0938052e-009 wkt1=-5.9083454e-008            pkt1=3.895127e-015              kt2=-0.067460028 ute=-1.8081944                 lute=3.1017917e-008             wute=3.3207417e-007 pute=-1.6935783e-014            ua1=4.451177e-010              lua1=-4.4203582e-018 wua1=2.7673753e-016             pua1=-1.8438104e-023            ub1=-1.1390928e-018 lub1=6.4971063e-026             wub1=1.6441283e-025             pub1=-6.5215153e-033 uc1=1.6354167e-013             luc1=8.0343594e-018             wuc1=8.6997706e-017 puc1=-3.1754592e-024            at=-3107.5194 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=2.3230473e-010             pcit=-1.285944e-017             lkt2=6.1251142e-010 lat=0.0030219345               wat=0.014394672                pat=-1.0570525e-009 letab=3.2438134e-008             petab=-2.7767585e-015            leta0=6.1625e-010 wkt2=-4.1887148e-009            pkt2=3.3871565e-018             u0_ff=-0.000304097 u0_ss=0.000483334                lu0_ff=1.5509e-11                 lu0_ss=-2.465e-11 wu0_ff=1.66037e-10                wu0_ss=3.3e-16                    pu0_ff=-8.46789e-18 pu0_ss=3.5e-23                    vsat_ff=-999.991                   vsat_ss=999.991 lvsat_ff=1.7e-10                    lvsat_ss=-1.7e-10                   wvsat_ff=1.7e-09 wvsat_ss=-1.7e-09                   pvsat_ff=1.7e-16                    pvsat_ss=-1.7e-16 a0_ff=0.241666                   a0_ss=-0.241666                  a0_sf=0.241666 la0_ff=-1.2325e-08                la0_ss=1.2325e-08                 la0_sf=-1.2325e-08 wa0_ff=1.7e-13                    wa0_ss=-1.7e-13                   wa0_sf=1.7e-13 pa0_ff=1.7e-20                    pa0_ss=-1.7e-20                   pa0_sf=1.7e-20 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.13 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.3589906 lvth0=-3.1637796e-009            wvth0=-2.2475401e-008            pvth0=1.2170775e-015 k2=0.042706517                lk2=-2.548934e-009             wk2=-1.0474856e-008 pk2=5.6125218e-016             cit=-0.00023237099             wcit=-5.480506e-009 voff=-0.085978835               lvoff=-5.8836216e-009            wvoff=-2.2724374e-008 pvoff=1.3584832e-015             eta0=0.14280978                 weta0=2.6675861e-008 etab=-0.51380191                wetab=8.4714193e-008             u0=0.0089845608 lu0=3.1893871e-010             wu0=6.6587571e-009             pu0=-2.8276758e-016 ua=-2.2405928e-009            lua=5.7565984e-017             wua=5.5255183e-016 pua=-2.208861e-023             ub=1.8021306e-018             lub=-4.3731785e-026 wub=-3.7120782e-025            pub=1.1873043e-032             uc=4.615227e-012 luc=-1.9733561e-018            wuc=1.6007265e-017             puc=-1.183886e-025 vsat=30276.232                  lvsat=0.0029846098               wvsat=0.021083967 pvsat=-9.1023201e-010            a0=-3.0612242                 la0=-2.3095739e-007 wa0=8.5435391e-006             pa0=-4.1361552e-013            ags=2 lags=0                          wags=0                          pags=0 keta=-0.20663617                lketa=5.8512725e-009             wketa=4.5947069e-008 pketa=-1.5197062e-015            pclm=0.20176053                 lpclm=4.6293158e-009 wpclm=1.2560465e-007             ppclm=-4.0022641e-015            pdiblc2=0.00033333333 lpdiblc2=2.38e-010                  wpdiblc2=0                          ppdiblc2=0 aigbacc=0.01579909                 laigbacc=-2.1206125e-010            waigbacc=-5.35136e-009 paigbacc=2.5534831e-016             aigc=0.0058107078               laigc=1.452618e-012 waigc=1.7914948e-010             paigc=-8.6496816e-018            aigsd=0.0056388035 laigsd=-2.3654547e-011            waigsd=-4.4327726e-010            paigsd=2.3264591e-017 tvoff=-0.00091126                ltvoff=9.72257e-011               wtvoff=2.13727e-009 ptvoff=-8.93197e-017              kt1=-0.28592369                lkt1=2.8227319e-009 wkt1=6.5170261e-008             pkt1=-2.4418125e-015            kt2=-0.069605551 ute=-1.2                       ua1=-5.5949557e-010            lua1=4.6814919e-017 wua1=1.1951235e-015             pua1=-6.5275787e-023            ub1=2.3851528e-018 lub1=-1.1476546e-025            wub1=-2.4327944e-024            pub1=1.2593605e-031 uc1=2.634e-010                 luc1=-5.3907e-018               wuc1=-3.29784e-017 puc1=2.9433222e-024             at=85651.568 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=1.6496238e-010             pcit=2.7855759e-016             lkt2=7.219331e-010 lat=-0.001504779               wat=-0.039786596               pat=1.7061921e-009 letab=2.0015501e-008             petab=-3.4327336e-015            leta0=1.1170133e-010 peta0=-1.3604689e-015            wkt2=8.7026333e-009             pkt2=-6.540716e-016 vsat_ff=-999.998                   vsat_ss=999.998                    lvsat_ff=6.7e-10 lvsat_ss=-6.7e-10                   wvsat_ff=-3.3e-09                   wvsat_ss=3.3e-09 pvsat_ff=2e-16                      pvsat_ss=-2e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.14 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.34026394 lvth0=-3.9502992e-009            wvth0=-3.8283357e-008            pvth0=1.8810116e-015 k2=0.008584745                lk2=-1.1158196e-009            wk2=-5.2269238e-009 pk2=3.4083903e-016             cit=-0.016311214               wcit=3.7183358e-009 voff=-0.096601918               lvoff=-5.4374521e-009            wvoff=-2.4424385e-008 pvoff=1.4298836e-015             eta0=0.12885689                 weta0=-2.6675861e-008 etab=-0.19223137                wetab=1.194663e-008              u0=0.017568415 lu0=-4.1583173e-011            wu0=-1.7291652e-009            pu0=6.9525158e-017 ua=-2.3774868e-009            lua=6.3315532e-017             wua=7.9805863e-016 pua=-3.2399895e-023            ub=3.4050451e-018             lub=-1.1105419e-025 wub=-1.6304665e-024            pub=6.4761908e-032             uc=2.8712827e-011 luc=-2.9854553e-018            wuc=2.2837193e-017             puc=-4.0524561e-025 vsat=94971.068                  lvsat=0.00026742667              wvsat=-0.0081789308 pvsat=3.1880971e-010             a0=33.385689                  la0=-1.7617277e-006 wa0=-6.0874309e-006            pa0=2.0088522e-013             ags=2 lags=0                          wags=0                          pags=0 keta=0.13259396                 lketa=-8.3963928e-009            wketa=-1.0386329e-008 pketa=8.462965e-016              pclm=0.48879756                 lpclm=-7.4262393e-009 wpclm=6.8906535e-008             ppclm=-1.6209433e-015            pdiblc2=-0.0068944444 lpdiblc2=5.4156667e-010             wpdiblc2=5.0383667e-009             ppdiblc2=-2.116114e-016 aigbacc=0.011183221                laigbacc=-1.8194745e-011            waigbacc=2.6785597e-009 paigbacc=-8.1908319e-017            aigc=0.0062269947               laigc=-1.6031434e-011 waigc=-2.5280763e-010            paigc=9.4925171e-018             aigsd=0.0045851903 laigsd=2.0597207e-011             waigsd=5.5495558e-010             paigsd=-1.8661188e-017 tvoff=0.000943991                ltvoff=1.93052e-011               wtvoff=9.09942e-010 ptvoff=-3.77721e-017              kt1=-0.33498695                lkt1=4.8833889e-009 wkt1=1.3636776e-007             pkt1=-5.4321074e-015            kt2=-0.089083338 ute=-1.7372033                 lute=2.256254e-008              wute=4.8670622e-007 pute=-2.0441661e-014            ua1=2.1034985e-009             lua1=-6.5030833e-017 wua1=1.3383692e-016             pua1=-2.0701752e-023            ub1=-2.7275257e-018 lub1=9.9967034e-026             wub1=3.0439644e-026             pub1=2.2480223e-032 uc1=3.501e-010                 luc1=-9.0321e-018               wuc1=-8.2446e-018 puc1=1.9045026e-024             at=53334.361 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=8.4027378e-010             pcit=-1.0779376e-016            lkt2=1.5400001e-009 lat=-0.0001474563              wat=-0.012518427               pat=5.6092907e-010 letab=6.5095384e-009             petab=-3.7649591e-016            leta0=6.9772267e-010 peta0=8.8030342e-016             wkt2=-6.8705e-009               pkt2=4.9715104e-029 vth0_ss=0.0184556                  vth0_mc=0.121611                   lvth0_ss=-7.75133e-10 lvth0_mc=-5.10767e-09               wvth0_ss=-1.00767e-08               wvth0_mc=-5.03837e-08 pvth0_ss=4.23223e-16                pvth0_mc=2.11612e-15                cit_mc=-0.01067 wcit_mc=3.02299e-09                voff_mc=0.0738222                  voff_mcl=0.0166833 lvoff_mc=-3.10053e-09               lvoff_mcl=-7.007e-10                 wvoff_mc=-4.03069e-08 wvoff_mcl=-1.51151e-08               pvoff_mc=1.69289e-15                pvoff_mcl=6.34834e-16 u0_ss=-0.00222444                u0_ff=0.00166833                 u0_sf=0.00278056 u0_mc=-0.000910554               lu0_ss=9.34267e-11                lu0_ff=-7.007e-11 lu0_sf=-1.16783e-10               lu0_mc=3.82437e-11                wu0_ss=2.01535e-09 wu0_ff=-1.51151e-09               wu0_sf=-2.51918e-09               wu0_mc=-5.03833e-10 pu0_ss=-8.46446e-17               pu0_ff=6.34834e-17                pu0_sf=1.05806e-16 pu0_mc=2.11611e-17                vsat_ff=-9445.52                   vsat_ss=773.882 vsat_sf=-4601.66                   vsat_fs=-11122.2                   vsat_mc=-31350 lvsat_ff=0.000354714                lvsat_ss=9.49667e-06                lvsat_sf=0.00019327 lvsat_fs=0.000467133                lvsat_mc=0.0013167                  wvsat_ff=0.00100768 wvsat_ss=0.00352686                 wvsat_sf=0.00151151                 wvsat_fs=0.0100767 wvsat_mc=0.0151151                  pvsat_ff=-4.23216e-11               pvsat_ss=-1.48128e-10 pvsat_sf=-6.34833e-11               pvsat_fs=-4.23223e-10               pvsat_mc=-6.34835e-10 lcit_mc=4.4814e-10                 pcit_mc=-1.26967e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.15 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.36657223 lvth0=-2.100185e-008             wvth0=-9.6035572e-009            pvth0=6.4557111e-015 k2=0.023766133                lk2=2.0058205e-013             wk2=2.1222751e-011 pk2=-1.2311776e-019            cit=0.0035088889               wcit=-2.2325333e-010 voff=-0.10752499                lvoff=-2.0816549e-008            wvoff=-4.9386497e-009 pvoff=3.5699547e-015             eta0=0.15022222                 weta0=-5.5813333e-009 etab=-0.32278778                wetab=6.2231867e-009             u0=0.014058885 lu0=0                          wu0=1.1689712e-010             pu0=0 ua=1.1857911e-009             lua=-3.6620508e-016            wua=-9.8410738e-017 pua=8.4683321e-023             ub=8.7680769e-019             lub=-6.0860198e-026 wub=-5.5555721e-026            pub=1.8809783e-032             uc=7.8366499e-011 luc=-3.3410415e-023            wuc=-8.8683495e-018            puc=1.3346099e-029 vsat=82146.719                  lvsat=4.684986e-008              wvsat=-0.0017185455 pvsat=-2.5580023e-014            a0=4.0106273                  la0=-1.515069e-006 wa0=-6.5136753e-007            pa0=4.1815906e-013             ags=1.47433 lags=1.2428114e-008             wags=-3.4243479e-007            pags=1.6956545e-013 keta=0.019777778                wketa=5.5813333e-009             pclm=0.26209243 lpclm=4.0963073e-012             wpclm=-6.6024687e-009            ppclm=-2.2365838e-018 pdiblc2=0.0011060812               lpdiblc2=-6.4171679e-010            wpdiblc2=-3.8662407e-011 ppdiblc2=1.7711381e-016             aigbacc=0.012781677                laigbacc=-1.0828028e-011 waigbacc=-2.370435e-010             paigbacc=2.9394227e-018             aigc=0.005998262 laigc=-3.6482818e-011            waigc=-1.1561961e-011            paigc=6.4564313e-018 aigsd=0.0048781314               laigsd=5.2223518e-011             waigsd=7.5257058e-011 paigsd=-2.8514035e-017            tvoff=0.000209892                ltvoff=6.66222e-010 wtvoff=1.14368e-010               ptvoff=-1.34718e-016              kt1=-0.26887876 lkt1=5.233809e-008              wkt1=1.6706281e-008             pkt1=-1.4321444e-014 kt2=-0.07                      ute=-1.1358275                 lute=-1.1203227e-013 wute=3.9873011e-008             pute=6.1169621e-020             ua1=2.1181187e-009 lua1=-5.1925972e-016            wua1=-9.1887469e-017            pua1=6.1753185e-023 ub1=-6.6376216e-019            lub1=-3.3820022e-025            wub1=3.8594623e-026 pub1=8.7627332e-032             uc1=3.5190837e-010             luc1=-1.2693301e-016 wuc1=1.1292898e-018             puc1=3.503351e-023              at=80000 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' a0_ff=-0.314534                  a0_ss=0.428063                   a0_sf=-0.303474 a0_fs=0.337872                   la0_ff=5.51238e-07                la0_ss=-6.53073e-07 la0_sf=4.51616e-07                la0_fs=-3.01077e-07               wa0_ff=9.29794e-08 wa0_ss=-1.54966e-07               wa0_sf=9.29796e-08                wa0_fs=-1.178e-07 pa0_ff=-8.34033e-14               pa0_ss=1.39005e-13                pa0_sf=-8.34032e-14 pa0_fs=5.56022e-14 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.16 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.37960699 lvth0=-9.3096661e-009            wvth0=-4.4165217e-009            pvth0=1.8029403e-015 k2=0.02329321                 lk2=4.2441244e-010             wk2=8.7438147e-010 pk2=-7.6540649e-016            cit=0.0051708283               wcit=-4.900366e-010 voff=-0.11702791                lvoff=-1.2292427e-008            wvoff=-2.3547199e-009 pvoff=1.2521697e-015             eta0=0.15022222                 weta0=-5.5813333e-009 etab=-0.32278778                wetab=6.2231867e-009             u0=0.013322118 lu0=6.6087941e-010             wu0=1.158016e-010              pu0=9.8268053e-019 ua=1.3021555e-009             lua=-4.7058398e-016            wua=-1.283295e-017 pua=7.9200456e-024             ub=6.2809276e-019             lub=1.6223709e-025 wub=-4.165376e-026             pub=6.3397242e-033             uc=6.2961909e-011 luc=1.3817884e-017             wuc=-1.1984583e-017            puc=2.7952751e-024 vsat=96997.761                  lvsat=-0.013321337               wvsat=-0.0098272142 pvsat=7.2734502e-009             a0=3.6928295                  la0=-1.2300043e-006 wa0=-5.1819744e-007            pa0=2.9870549e-013             ags=2.08477 lags=-5.3513653e-007            wags=-3.3873907e-007            pags=1.6625039e-013 keta=0.019998518                lketa=-1.9800444e-010            wketa=3.7208889e-011 pketa=4.9730796e-015             pclm=0.26808742                 lpclm=-5.3734108e-009 wpclm=-6.875572e-009             ppclm=2.4273701e-016             pdiblc2=-0.0012810248 lpdiblc2=1.4995173e-009             wpdiblc2=3.5643687e-010             ppdiblc2=-1.7729025e-016 aigbacc=0.013746671                laigbacc=-8.7642745e-010            waigbacc=-4.0880682e-010 paigbacc=1.5701111e-016             aigc=0.0059530337               laigc=4.0869424e-012 waigc=-4.1672289e-012            paigc=-1.7664379e-019            aigsd=0.004936492 laigsd=-1.2598449e-013            waigsd=4.3392155e-011             paigsd=6.8782664e-020 tvoff=0.000238657                ltvoff=6.40419e-010               wtvoff=1.46741e-010 ptvoff=-1.63756e-016              kt1=-0.24474059                lkt1=3.0686156e-008 wkt1=9.6674403e-009             pkt1=-8.0076041e-015            kt2=-0.07 ute=-1.2586951                 lute=1.102121e-007              wute=1.3098525e-007 pute=-8.172762e-014             ua1=2.0962901e-009             lua1=-4.9967946e-016 wua1=-9.4507369e-017            pua1=6.4103235e-023             ub1=-1.2862835e-018 lub1=2.2020141e-025             wub1=3.615246e-025              pub1=-2.0204086e-031 uc1=-4.8572242e-011            luc1=2.322981e-016              wuc1=1.1659682e-016 puc1=-6.8540863e-023            at=70066.667 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=-1.4907596e-009            pcit=2.3930459e-016             lat=0.0089102 u0_ff=0.000149                   u0_ss=-9.93333e-05               u0_sf=4.85629e-05 u0_fs=-9.93333e-05               lu0_ff=-1.33653e-10               lu0_ss=8.9102e-11 lu0_sf=-4.35609e-11               lu0_fs=8.9102e-11                 wu0_ff=-3.3e-17 wu0_ss=-4.4e-17                   wu0_sf=2.77207e-11                wu0_fs=-4.4e-17 pu0_ff=6e-24                      pu0_ss=-4e-24                     pu0_sf=-2.48654e-17 pu0_fs=-4e-24                     a0_ff=0.300001                   a0_ss=-0.300001 a0_sf=0.200001                   a0_fs=0.0423975                  la0_ff=-1.3e-13 la0_ss=1.3e-13                    la0_sf=-9e-14                     la0_fs=-3.60369e-08 wa0_ff=2.7e-13                    wa0_ss=-2.7e-13                   wa0_sf=-4.9e-13 wa0_fs=-6.69015e-08               pa0_ff=-6.1e-19                   pa0_ss=6.1e-19 pa0_sf=-7e-21                     pa0_fs=9.94641e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.17 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.39962082 lvth0=-3.6348695e-010            wvth0=5.5106844e-011             pvth0=-1.9587768e-016 k2=0.019717986                lk2=2.0225378e-009             wk2=4.0548812e-010 pk2=-5.5581116e-016            cit=0.00025141143              wcit=4.1559845e-010 voff=-0.14097156                lvoff=-1.5896194e-009            wvoff=3.8516308e-010 pvoff=2.7442037e-017             eta0=0.15022222                 weta0=-5.5813333e-009 etab=-0.32278778                wetab=6.2231867e-009             u0=0.013491697 lu0=5.8507773e-010             wu0=1.6653805e-010             pu0=-2.1696512e-017 ua=1.0565394e-009             lua=-3.607936e-016             wua=8.3563809e-018 pua=-1.5515855e-024            ub=8.3369591e-019             lub=7.0332479e-026 wub=-6.4692498e-026            pub=1.663804e-032              uc=8.6849251e-011 luc=3.1402421e-018             wuc=-1.2898512e-017            puc=3.2038013e-024 vsat=53334.977                  lvsat=0.0061959268               wvsat=0.014254523 pvsat=-3.4910864e-009            a0=2.0197113                  la0=-4.8212052e-007 wa0=2.6947853e-007             pa0=-5.3385669e-014            ags=-0.58010405 lags=6.5606216e-007             wags=6.3393296e-008             pags=-1.3502772e-014 keta=0.095921011                lketa=-3.4135359e-008            wketa=-7.1287222e-010 pketa=5.3083659e-015             pclm=0.082252446                lpclm=7.7694825e-008 wpclm=2.1533205e-009             ppclm=-3.793178e-015             pdiblc2=0.0012303385 lpdiblc2=3.7693791e-010             wpdiblc2=-7.67648e-011              ppdiblc2=1.6350902e-017 aigbacc=0.012635835                laigbacc=-3.7988384e-010            waigbacc=-5.1327857e-010 paigbacc=2.0370999e-016             aigc=0.005932246                laigc=1.337903e-011 waigc=7.2817468e-012             paigc=-5.2943359e-018            aigsd=0.0049121966 laigsd=1.0734089e-011             waigsd=3.7892076e-011             paigsd=2.5273181e-018 tvoff=0.00204062                 ltvoff=-1.65059e-010              wtvoff=-3.8685e-010 ptvoff=7.4759e-017                kt1=-0.1405518                 lkt1=-1.5886236e-008 wkt1=-1.6675208e-008            pkt1=3.7675597e-015             kt2=-0.07 ute=-0.84113056                lute=-7.6439234e-008            wute=-9.9047966e-008 pute=2.1097229e-014             ua1=1.0658274e-009             lua1=-3.9062641e-017 wua1=5.7344137e-017             pua1=-3.7743878e-024            ub1=-1.2031627e-018 lub1=1.8304643e-025             wub1=-9.5181324e-026            pub1=2.1066911e-033 uc1=6.5799534e-010             luc1=-8.3537607e-017            wuc1=-7.4752251e-017 puc1=1.6992171e-023             at=135710.54 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=7.082197e-010              pcit=-1.6551428e-016            lat=-0.020432609 wat=-0.0038327798              pat=1.7132526e-009             u0_ff=-5.8974e-05 u0_ss=5.44873e-05                u0_sf=4.2137e-05                 u0_fs=5.44873e-05 lu0_ff=-4.06887e-11               lu0_ss=2.03446e-11                lu0_sf=-4.06883e-11 lu0_fs=2.03446e-11                wu0_ff=3.3e-16                    wu0_ss=-2.2e-16 wu0_sf=-2.79067e-11               wu0_fs=-2.2e-16                   pu0_ff=-2e-23 pu0_ss=1.3e-23                    pu0_sf=-2e-23                     pu0_fs=1.3e-23 a0_ff=0.254489                   a0_ss=-0.300001                  a0_sf=0.200001 a0_fs=-0.0750379                 la0_ff=2.03447e-08                la0_ss=-5e-14 la0_sf=2.01e-13                   la0_fs=1.64562e-08                wa0_ff=4.4e-13 wa0_ss=3.3e-13                    wa0_sf=1.1e-13                    wa0_fs=-3.44901e-08 pa0_ff=-4.7e-20                   pa0_ss=-6e-20                     pa0_sf=7.3e-20 pa0_fs=-4.54187e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.18 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.3919791 lvth0=-1.9911737e-009            wvth0=-3.7195117e-009            pvth0=6.0811606e-016 k2=0.043035032                lk2=-2.9439931e-009            wk2=-5.2279105e-009 pk2=6.4410274e-016             cit=0.0054543758               wcit=-7.6857928e-010 voff=-0.13019769                lvoff=-3.8844519e-009            wvoff=-1.9038027e-009 pvoff=5.1499174e-016             eta0=0.15022222                 weta0=-5.5813333e-009 etab=-0.32278498                wetab=6.2214679e-009             u0=0.015939283 lu0=6.3742002e-011             wu0=-1.6614712e-011            pu0=1.7315026e-017 ua=-3.9498309e-010            lua=-5.1619303e-017            wua=5.7853604e-018 pua=-1.0039581e-024            ub=1.3334886e-018             lub=-3.6123363e-026 wub=2.6836794e-026             pub=-2.8576991e-033            uc=1.5223707e-010 luc=-1.0787363e-017            wuc=5.5142139e-018             puc=-7.1810937e-025 vsat=92805.429                  lvsat=-0.0022112795              wvsat=-0.0087479386 pvsat=1.408438e-009              a0=2.8392763                  la0=-6.5668787e-007 wa0=-4.6098994e-007            pa0=1.0220412e-013             ags=2.8452381 lags=-7.3535714e-008            wags=0                          pags=0 keta=-0.053064947               lketa=-2.4013496e-009            wketa=2.9363461e-008 pketa=-1.0978931e-015            pclm=0.47673865                 lpclm=-6.3307368e-009 wpclm=-2.6129901e-008            ppclm=2.2311482e-015             pdiblc2=0.0023095238 lpdiblc2=1.4707143e-010             wpdiblc2=0                          ppdiblc2=0 aigbacc=0.011432988                laigbacc=-1.2367746e-010            waigbacc=4.4375294e-010 paigbacc=-1.37723e-019              aigc=0.0060257027               laigc=-6.5272358e-012 waigc=-2.2976312e-011            paigc=1.1506306e-018             aigsd=0.0048835312 laigsd=1.6839802e-011             waigsd=5.4968559e-011             paigsd=-1.1099728e-018 tvoff=0.00147578                 ltvoff=-4.47481e-011              wtvoff=-9.32111e-011 ptvoff=1.22139e-017               kt1=-0.2251901                 lkt1=2.1417231e-009 wkt1=4.2656477e-009             pkt1=-6.9284255e-016            kt2=-0.0723011 ute=-1.1294183                 lute=-1.5033938e-008            wute=-3.8537683e-008 pute=8.2085385e-015             ua1=1.1403439e-009             lua1=-5.4934657e-017 wua1=6.5441924e-017             pua1=-5.4992164e-024            ub1=-2.5082905e-019 lub1=-1.9800643e-026            wub1=-2.384157e-025             pub1=3.2615613e-032 uc1=3.47e-010                  luc1=-1.72956e-017              wuc1=-5.382e-018 puc1=2.2163076e-024             at=45277.3                    jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)' jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 lcit=-4.0001171e-010 pcit=8.6715579e-017             lkt2=4.9013435e-010             lat=-0.0011703302 wat=0.0056427436               pat=-3.050339e-010             letab=-5.9550856e-013 petab=3.6610118e-019             wkt2=5.0994074e-010             pkt2=-1.0861738e-016 u0_ff=-0.000422619               u0_ss=0.000115477                u0_sf=-0.000251693 u0_fs=0.000253572                lu0_ff=3.67679e-11                lu0_ss=7.35355e-12 lu0_sf=2.18973e-11                lu0_fs=-2.20607e-11               wu0_ff=2.2e-16 wu0_ss=-3.3e-16                   wu0_sf=-4.71758e-11               wu0_fs=-3.3e-16 pu0_ff=-3.3e-23                   pu0_ss=-2e-23                     pu0_sf=4.10427e-18 pu0_fs=-2e-23                     vsat_ff=690.48                     vsat_ss=-690.48 lvsat_ff=-0.000147071               lvsat_ss=0.000147071                wvsat_ff=-2.2e-10 wvsat_ss=2.2e-10                    pvsat_ff=3.3e-17                    pvsat_ss=-3.3e-17 a0_ff=0.522617                   a0_ss=-0.438099                  a0_sf=0.198466 a0_fs=0.00375647                 la0_ff=-3.6768e-08                la0_ss=2.94143e-08 la0_sf=3.26837e-10                la0_fs=-3.26837e-10               wa0_ff=1.22e-13 wa0_ss=-5.22e-13                  wa0_sf=3.85382e-08                wa0_fs=-9.43511e-08 pa0_ff=3.67e-20                   pa0_ss=-6.7e-21                   pa0_sf=-8.20854e-15 pa0_fs=8.20854e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.19 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.40315175 lvth0=-1.0191527e-009            wvth0=4.3039285e-009             pvth0=-8.9923233e-017 k2=0.042165868                lk2=-2.8683758e-009            wk2=-7.563927e-010 pk2=2.5508069e-016             cit=-0.002909665               wcit=9.7439671e-010 voff=-0.1347819                 lvoff=-3.4856262e-009            wvoff=2.7821182e-009 pvoff=1.0731663e-016             eta0=0.13589815                 weta0=-1.6278889e-009 etab=-0.63436482                wetab=4.6840407e-009             u0=0.015446472 lu0=1.0661657e-010             wu0=6.4030521e-010             pu0=-3.9837007e-017 ua=-1.0749028e-009            lua=7.5337105e-018             wua=-4.0277317e-017 pua=3.0034948e-024             ub=1.1406931e-018             lub=-1.9350154e-026 wub=3.9712191e-026             pub=-3.9778586e-033            uc=7.3686429e-011 luc=-3.9534573e-018            wuc=-2.6148125e-018            puc=-1.0884081e-026 vsat=30067.912                  lvsat=0.0032468845               wvsat=0.017214393 pvsat=-8.5028486e-010            a0=-3.5671258                 la0=-9.9330879e-008 wa0=2.7159376e-006             pa0=-1.7418858e-013            ags=2 lags=0                          wags=0                          pags=0 keta=-0.16060368                lketa=6.9545205e-009             wketa=6.9925767e-008 pketa=-4.6268137e-015            pclm=0.41334449                 lpclm=-8.1544509e-010 wpclm=1.3144486e-008             ppclm=-1.1857234e-015            pdiblc2=0.0025833333 lpdiblc2=1.2325e-010                wpdiblc2=0                          ppdiblc2=0 aigbacc=0.010188225                laigbacc=-1.5383017e-011            waigbacc=1.9961076e-010 paigbacc=2.1102647e-017             aigc=0.0060217737               laigc=-6.1854141e-012 waigc=1.0325701e-011             paigc=-1.7466445e-018            aigsd=0.0050223152 laigsd=4.7656025e-012             waigsd=3.7930774e-011             paigsd=3.7231451e-019 tvoff=-0.000284382               ltvoff=1.08386e-010               wtvoff=2.2148e-010 ptvoff=-1.51642e-017              kt1=-0.21247997                lkt1=1.0359415e-009 wkt1=-3.724328e-009             pkt1=2.2853392e-018             kt2=-0.067518371 ute=-1.2807896                 lute=-1.8646356e-009            wute=4.4111138e-008 pute=1.018091e-015              ua1=9.1230091e-010             lua1=-3.5094913e-017 wua1=2.1655493e-017             pua1=-1.6897969e-024            ub1=-9.6960701e-019 lub1=4.273304e-026              wub1=7.1873584e-026             pub1=5.6204453e-033 uc1=8.36e-011                  luc1=5.6202e-018                wuc1=4.14414e-017 puc1=-1.8573282e-024            at=10651.021 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=3.2765984e-010             pcit=-6.4923332e-017            lkt2=7.4036938e-011 lat=0.001842156                wat=0.0068825086               pat=-4.1289346e-010 letab=2.710685e-008              petab=1.3412226e-016             leta0=1.2461944e-009 peta0=-3.4394967e-016            wkt2=-4.1568592e-009            pkt2=2.9739422e-016 u0_ss=0.000483333                lu0_ss=-2.465e-11                 wu0_ss=4.4e-16 pu0_ss=1.3e-23                    vsat_ff=448.14                     vsat_ss=1000.01 lvsat_ff=-0.000125989               lvsat_ss=1.1e-10                    wvsat_ff=-0.000790691 wvsat_ss=2.11e-09                   pvsat_ff=6.879e-11                  pvsat_ss=-6.7e-17 a0_ff=0.241667                   a0_ss=-0.241667                  a0_sf=0.488704 la0_ff=-1.2325e-08                la0_ss=1.2325e-08                 la0_sf=-2.49239e-08 wa0_ff=2.2e-13                    wa0_ss=-2.2e-13                   wa0_sf=-1.34882e-07 pa0_ff=-3.3e-21                   pa0_ss=3.3e-21                    pa0_sf=6.87899e-15 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.20 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.41862252 lvth0=-2.3014367e-010            wvth0=1.0083625e-008             pvth0=-3.8468777e-016 k2=0.020482556                lk2=-1.7625269e-009            wk2=1.6594264e-009 pk2=1.3187392e-016             cit=-0.017211768               wcit=3.790245e-009 voff=-0.14538816                lvoff=-2.9447069e-009            wvoff=9.7131163e-009 pvoff=-2.4616427e-016            eta0=0.23085185                 weta0=-2.1395111e-008 etab=-0.40737364                wetab=2.6604355e-008             u0=0.022356897 lu0=-2.4581512e-010            wu0=-6.4253835e-010            pu0=2.5588014e-017 ua=-1.3468646e-009            lua=2.1403761e-017             wua=6.4576235e-017 pua=-2.3440363e-024            ub=1.4204298e-018             lub=-3.3616728e-026 wub=-1.6279918e-025            pub=6.3502211e-033             uc=2.8104537e-011 luc=-1.6287808e-018            wuc=3.1821015e-018             puc=-3.0652669e-025 vsat=94595.629                  lvsat=-4.402903e-005             wvsat=-0.014034424 pvsat=7.4340478e-010             a0=25.138133                  la0=-1.5632991e-006 wa0=-6.8533102e-006            pa0=3.1384306e-013             ags=2 lags=0                          wags=0                          pags=0 keta=0.041533043                lketa=-3.3544526e-009            wketa=-8.9553319e-008 pketa=3.5066197e-015             pclm=0.45319897                 lpclm=-2.8480232e-009 wpclm=-1.1680737e-008            ppclm=8.0362962e-017             pdiblc2=0.00033333333 lpdiblc2=2.38e-010                  wpdiblc2=0                          ppdiblc2=0 aigbacc=-0.004632632               laigbacc=7.4048068e-010             waigbacc=5.8043604e-009 paigbacc=-2.6473958e-016            aigc=0.0062698406               laigc=-1.8836825e-011 waigc=-7.1537017e-011            paigc=2.4283541e-018             aigsd=0.0045139546 laigsd=3.0691993e-011             waigsd=1.7089028e-010             paigsd=-6.4086201e-018 tvoff=0.00489467                 ltvoff=-1.55745e-010              wtvoff=-1.03277e-009 ptvoff=4.88025e-017               kt1=-0.10017476                lkt1=-4.6916244e-009 wkt1=-3.6248657e-008            pkt1=1.6610261e-015             kt2=-0.047192583 ute=-1.3879526                 lute=3.6006756e-009             wute=1.0262212e-007 pute=-1.9659689e-015            ua1=1.7005049e-009             lua1=-7.5293318e-017 wua1=-3.8836805e-017            pua1=1.3953103e-024             ub1=-3.1648404e-018 lub1=1.5468994e-025             wub1=5.975019e-025              pub1=-2.1186599e-032 uc1=1.5086667e-010             luc1=2.1896e-018                wuc1=2.84648e-017 puc1=-1.1955216e-024            at=15710.866 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=1.0570671e-009             pcit=-2.0853159e-016            lkt2=-9.6257826e-010 lat=0.0015841039               wat=-0.0015989725              pat=1.966208e-011 letab=1.55303e-008               petab=-9.8381376e-016            leta0=-3.5964444e-009 peta0=6.6417867e-016             wkt2=-3.534847e-009             pkt2=2.656716e-016 vsat_ff=-6792.63                   vsat_ss=1000.04                    lvsat_ff=0.000243289 lvsat_ss=1.1e-10                    wvsat_ff=0.00316276                 wvsat_ss=-2.2e-09 pvsat_ff=-1.32836e-10               pvsat_ss=7.3e-16 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.21 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=2.7e-007                   wmax=5.4e-007                   vth0=-0.42183778 lvth0=-9.510256e-011             wvth0=6.2559588e-009             pvth0=-2.2392577e-016 k2=-0.0020439242              lk2=-8.1641472e-010            wk2=5.7632958e-010 pk2=1.7736399e-016             cit=-0.0014689604              wcit=-4.3855345e-009 voff=-0.14531384                lvoff=-2.9478281e-009            wvoff=2.1723266e-009 pvoff=7.0548894e-017             eta0=0.052740741                weta0=1.4883556e-008 etab=-0.19994609                wetab=1.6158865e-008             u0=0.015810505 lu0=2.9133333e-011             wu0=-7.6934624e-010            pu0=3.0913946e-017 ua=-8.8193885e-010            lua=1.8768814e-018             wua=-1.8510528e-017 pua=1.1456077e-024             ub=3.8472688e-019             lub=9.8827961e-027 wub=1.8627227e-026             pub=-1.2696878e-033            uc=1.4409159e-010 luc=-6.5002369e-018            wuc=-4.015961e-017             puc=1.5138252e-024 vsat=68853.192                  lvsat=0.0010371533               wvsat=0.0060814292 pvsat=-1.0146104e-010            a0=32.550844                  la0=-1.874633e-006 wa0=-5.6316061e-006            pa0=2.6253148e-013             ags=2 lags=0                          wags=0                          pags=0 keta=0.28221628                 lketa=-1.3463149e-008            wketa=-9.2080116e-008 pketa=3.6127452e-015             pclm=0.98813837                 lpclm=-2.5315478e-008 wpclm=-2.0373355e-007            ppclm=8.1465811e-015             pdiblc2=-0.005162963 lpdiblc2=4.6884444e-010             wpdiblc2=4.0929778e-009             ppdiblc2=-1.7190507e-016 aigbacc=0.01914486                 laigbacc=-2.5817398e-010            waigbacc=-1.668495e-009 paigbacc=4.9120343e-017             aigc=0.0056319428               laigc=7.9548797e-012 waigc=7.2090708e-011             paigc=-3.6040103e-018            aigsd=0.0056020776 laigsd=-1.5009175e-011            waigsd=-2.6487706e-013            paigsd=7.7989633e-019 tvoff=0.000440132                ltvoff=3.13451e-011               wtvoff=1.18505e-009 ptvoff=-4.43459e-017              kt1=-0.15148149                lkt1=-2.5367414e-009 wkt1=3.617378e-008              pkt1=-1.3807162e-015            kt2=-0.1067778 ute=-0.32470518                lute=-4.1055716e-008            wute=-2.8451777e-007 pute=1.4293906e-014             ua1=3.5411637e-009             lua1=-1.5260099e-016 wua1=-6.5112827e-016            pua1=2.7111552e-023             ub1=-3.2349182e-018 lub1=1.5763321e-025             wub1=3.0747595e-025             pub1=-9.0055089e-033 uc1=2.338e-010                 luc1=-1.2936e-018               wuc1=5.52552e-017 puc1=-2.3207184e-024            at=56501.005 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=3.9586918e-010             pcit=1.3485115e-016             lkt2=1.5400006e-009 lat=-0.0001290819              wat=-0.014247415               pat=5.5089665e-010 letab=6.818343e-009              petab=-5.451032e-016             leta0=3.8842222e-009 peta0=-8.5952533e-016            wkt2=2.7906734e-009             pkt2=-2.578576e-022 vth0_mc=0.0293333                  lvth0_mc=-1.232e-09                 wvth0_mc=1.1e-14 pvth0_mc=-2.7e-22                   cit_mc=-0.0103807                 wcit_mc=2.86508e-09 voff_mcl=-0.0166222                 lvoff_mcl=6.98134e-10                wvoff_mcl=3.06974e-09 pvoff_mcl=-1.28929e-16               u0_ss=0.00296593                 u0_ff=-0.00222444 u0_sf=-0.00370741                u0_mc=-0.00370741                lu0_ss=-1.24569e-10 lu0_ff=9.34267e-11                lu0_sf=1.55711e-10                lu0_mc=1.55711e-10 wu0_ss=-8.18596e-10               wu0_ff=6.13947e-10                wu0_sf=1.02324e-09 wu0_mc=1.02324e-09                pu0_ss=3.4381e-17                 pu0_ff=-2.57858e-17 pu0_sf=-4.29763e-17               pu0_mc=-4.29763e-17               vsat_ss=9857.03 vsat_ff=-10598.5                   vsat_sf=-3707.41                   vsat_fs=1711.08 vsat_mc=81.4863                    vsat_mcl=7496.3                     lvsat_ss=-0.000371996 lvsat_ff=0.000403138                lvsat_sf=0.000155711                lvsat_fs=-7.18662e-05 lvsat_mc=-3.42244e-06               lvsat_mcl=-0.000314844               wvsat_ss=-0.00143254 wvsat_ff=0.00163719                 wvsat_sf=0.00102324                 wvsat_fs=0.00306973 wvsat_mc=-0.00204649                wvsat_mcl=-0.00409298                pvsat_ss=6.01665e-11 pvsat_ff=-6.87625e-11               pvsat_sf=-4.29763e-11               pvsat_fs=-1.28929e-10 pvsat_mc=8.59526e-11                pvsat_mcl=1.71905e-10                lcit_mc=4.35991e-10 pcit_mc=-1.20334e-16 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.22 pmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.38238507 lvth0=-9.1586792e-009            wvth0=-5.2392142e-009            pvth0=3.1869961e-015 k2=0.013545008                lk2=-7.1197321e-014            wk2=2.8422533e-009 pk2=-4.8106658e-020            cit=0.0024888889               wcit=5.8266667e-011 voff=-0.11962078                lvoff=-2.0047877e-008            wvoff=-1.6002125e-009 pvoff=3.3578014e-015             eta0=0.13576333                 weta0=-1.59068e-009 etab=-0.33207556                wetab=8.7866133e-009             u0=0.013801549 lu0=-9.3950648e-014            wu0=1.8792168e-010             pu0=2.5930379e-020 ua=9.2374155e-010             lua=-2.2379178e-016            wua=-2.6085076e-017 pua=4.5377251e-023             ub=7.9735982e-019             lub=-4.4127602e-027 wub=-3.362811e-026             pub=3.2302901e-033             uc=6.419001e-011 luc=1.0037147e-023             wuc=-4.9556384e-018            puc=1.354572e-030 vsat=57849.068                  lvsat=-7.80831e-008              wvsat=0.0049876063 pvsat=8.9014733e-015             a0=1.5933185                  la0=1.6974587e-013 wa0=1.5809691e-008             pa0=-1.9351029e-020            ags=0.13787064 lags=7.2134573e-007             wags=2.6428001e-008             pags=-2.6095806e-014 keta=0.061111111                wketa=-5.8266667e-009            pclm=0.23118998 lpclm=-6.5186842e-012            wpclm=1.9266074e-009             ppclm=6.9315386e-019 pdiblc2=0.00080133335              lpdiblc2=-1.4767891e-016            wpdiblc2=4.5447998e-011 ppdiblc2=1.6835395e-023             aigbacc=0.012064088                laigbacc=2.9983578e-012 waigbacc=-3.8988734e-011            paigbacc=-8.7665967e-019            aigc=0.0059752141 laigc=-3.3024624e-011            waigc=-5.2007524e-012            paigc=5.5019697e-018 aigsd=0.0051197554               laigsd=-1.0806799e-010            waigsd=8.5688207e-012 paigsd=1.5726421e-017             tvoff=0.000112084                ltvoff=6.49819e-010 wtvoff=1.41363e-010               ptvoff=-1.30191e-016              kt1=-0.22014254 lkt1=1.685925e-008              wkt1=3.2550838e-009             pkt1=-4.5292846e-015 kt2=-0.071116074               ute=-0.91490974                lute=1.8672045e-013 wute=-2.110029e-008             pute=-2.1286132e-020            ua1=2.2084699e-009 lua1=-6.0670576e-016            wua1=-1.1682439e-016            pua1=8.5888294e-023 ub1=-4.8187203e-019            lub1=3.1027997e-026             wub1=-1.1607052e-026 pub1=-1.4279655e-032            uc1=3.060558e-010              luc1=5.0480945e-017 wuc1=1.3784598e-017             puc1=-1.3932741e-023            at=80000 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' wkt2=3.0803644e-010             a0_ff=-0.157469                  a0_ss=0.011223 a0_sf=-0.115114                  a0_fs=-0.0576464                 la0_ff=2.84105e-07 la0_ss=-1.84483e-07               la0_sf=2.19537e-07                la0_fs=-6.45696e-08 wa0_ff=4.96296e-08                wa0_ss=-3.99185e-08               wa0_sf=4.09927e-08 wa0_fs=-8.63706e-09               pa0_ff=-9.67475e-15               pa0_ss=9.67437e-15 pa0_sf=-1.93487e-14               pa0_fs=-9.67435e-15               pdiblc2_sf=7.03704e-05 pdiblc2_fs=-7.03704e-05               lpdiblc2_sf=-5e-18                     lpdiblc2_fs=5e-18 wpdiblc2_sf=-1.94222e-11               wpdiblc2_fs=1.94222e-11                ppdiblc2_sf=-5e-23 ppdiblc2_fs=5e-23 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.23 pmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.38807586 lvth0=-4.0540336e-009            wvth0=-2.0791135e-009            pvth0=3.5238574e-016 k2=0.018803797                lk2=-4.7172051e-009            wk2=2.1134595e-009 pk2=6.5367994e-016             cit=0.0029745185               wcit=1.1614489e-010 voff=-0.13148878                lvoff=-9.4022782e-009            wvoff=1.6364796e-009 pvoff=4.5448854e-016             eta0=0.13576333                 weta0=-1.59068e-009 etab=-0.33207556                wetab=8.7866133e-009             u0=0.012750619 lu0=9.4259082e-010             wu0=2.735355e-010              pu0=-7.6769667e-017 ua=1.1991357e-009             lua=-4.7082031e-016            wua=1.5600518e-017 pua=7.985273e-024              ub=7.6648068e-019             lub=2.3285831e-026 wub=-7.9848824e-026            pub=4.4690271e-032             uc=7.1194658e-011 luc=-6.2831593e-018            wuc=-1.4256822e-017            puc=8.343163e-024 vsat=15797.537                  lvsat=0.037720145                wvsat=0.012584048 pvsat=-6.813999e-009             a0=1.5104798                  la0=7.4306466e-008 wa0=8.4131064e-008             pa0=-6.1284291e-014            ags=0.73141771 lags=1.8893401e-007             wags=3.4786158e-008             pags=-3.3593073e-014 keta=0.034254321                lketa=2.4090541e-008             wketa=-3.8973926e-009 pketa=-1.7305588e-015            pclm=0.21571442                 lpclm=1.3875064e-008 wpclm=7.579378e-009              ppclm=-5.0698421e-015            pdiblc2=-0.00030663832 lpdiblc2=9.9385044e-010             wpdiblc2=8.7506208e-011             ppdiblc2=-3.7726198e-017 aigbacc=0.012632718                laigbacc=-5.0706286e-010            waigbacc=-1.0135568e-010 paigbacc=5.5066486e-017             aigc=0.0059190583               laigc=1.734711e-011 waigc=5.2099718e-012             paigc=-3.8364499e-018            aigsd=0.005011627 laigsd=-1.1076805e-011            waigsd=2.2654898e-011             paigsd=3.091209e-018 tvoff=0.00112337                 ltvoff=-2.57306e-010              wtvoff=-9.74402e-011 ptvoff=8.4016e-017                kt1=-0.18745252                lkt1=-1.2463698e-008 wkt1=-6.1440693e-009            pkt1=3.9017557e-015             kt2=-0.072224708 ute=-0.63171966                lute=-2.5402131e-007            wute=-4.2059959e-008 pute=1.8800802e-014             ua1=1.7597935e-009             lua1=-2.0424305e-016 wua1=-1.6343057e-018            pua1=-1.7437213e-023            ub1=1.2977273e-019 lub1=-5.1761736e-025            wub1=-2.9306915e-026            pub1=1.5971227e-033 uc1=4.3683333e-010             luc1=-6.68265e-017              wuc1=-1.737512e-017 puc1=1.4017527e-023             at=70066.667                  pat=0 wat=0                          jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)' jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 lcit=-4.3560978e-010 pcit=-5.1916765e-017            lkt2=9.9444432e-010             lat=0.0089102 wkt2=6.1401931e-010             pkt2=-2.7446663e-016            u0_ff=9.19768e-06 u0_ss=-2.94325e-05               u0_sf=9.19768e-06                u0_fs=-2.94325e-05 lu0_ff=-8.25007e-12               lu0_ss=2.64002e-11                lu0_sf=-8.25007e-12 lu0_fs=2.64002e-11                wu0_ff=3.85855e-11                wu0_ss=-1.92928e-11 wu0_sf=3.85855e-11                wu0_fs=-1.92928e-11               pu0_ff=-3.46112e-17 pu0_ss=1.73056e-17                pu0_sf=-3.46112e-17               pu0_fs=1.73056e-17 vsat_mc=1398.02                    lvsat_mc=-0.00125403                wvsat_mc=-0.000385855 pvsat_mc=3.46112e-10                a0_ff=0.124304                   a0_ss=-0.159489 a0_sf=0.0597287                  a0_fs=-0.0597287                 la0_ff=3.13507e-08 la0_ss=-3.13514e-08               la0_sf=6.27012e-08                la0_fs=-6.27012e-08 wa0_ff=4.84907e-08                wa0_ss=-3.878e-08                 wa0_sf=3.8715e-08 wa0_fs=-3.8715e-08                pa0_ff=-8.65275e-15               pa0_ss=8.65275e-15 pa0_sf=-1.73055e-14               pa0_fs=1.73055e-14                pdiblc2_sf=0.000140272 pdiblc2_fs=-0.000140272               lpdiblc2_sf=-6.27014e-11               lpdiblc2_fs=6.27014e-11 wpdiblc2_sf=-3.8715e-11                wpdiblc2_fs=3.8715e-11                 ppdiblc2_sf=1.73056e-17 ppdiblc2_fs=-1.73056e-17               at_mc=-6291.11                   pat_mc=-1.5575e-09 wat_mc=0.00173635                 lat_mc=0.00564313 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.24 pmos ( level=54                         lmin=2.16e-007                  lmax=4.5e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.38999377 lvth0=-3.1967305e-009            wvth0=-2.6019587e-009            pvth0=5.8609753e-016 k2=0.005324174                lk2=1.3081865e-009             wk2=4.3781802e-009 pk2=-3.5865019e-016            cit=0.0019017074               wcit=-3.9883234e-011 voff=-0.14747857                lvoff=-2.2548408e-009            wvoff=2.1811002e-009 pvoff=2.1104313e-016             eta0=0.13576333                 weta0=-1.59068e-009 etab=-0.33207556                wetab=8.7866133e-009             u0=0.013527706 lu0=5.9523298e-010             wu0=1.5659969e-010             pu0=-2.4499359e-017 ua=8.4874729e-010             lua=-3.141967e-016             wua=6.570701e-017 pua=-1.4412329e-023            ub=6.7758888e-019             lub=6.3020461e-026 wub=-2.1606958e-026            pub=1.8656157e-032             uc=2.9856467e-012 luc=2.4206269e-017             wuc=1.0247843e-017             puc=-2.6104221e-024 vsat=121670.12                  lvsat=-0.0096048989              wvsat=-0.0046059758 pvsat=8.699415e-010              a0=3.8820915                  la0=-9.8580397e-007 wa0=-2.4453841e-007            pa0=8.5630963e-014             ags=-0.95653281 lags=9.4344789e-007             wags=1.6728763e-007             pags=-9.2821232e-014 keta=0.14494646                 lketa=-2.5388846e-008            wketa=-1.4243897e-008 pketa=2.8943285e-015             pclm=0.099251992                lpclm=6.5933768e-008 wpclm=-2.538554e-009             ppclm=-5.4712647e-016            pdiblc2=0.0022117987 lpdiblc2=-1.3189089e-010            wpdiblc2=-3.4764782e-010            ppdiblc2=1.5678765e-016 aigbacc=0.0098785416               laigbacc=7.2405387e-010             waigbacc=2.4773449e-010 paigbacc=-1.0097682e-016            aigc=0.0059685479               laigc=-4.7747424e-012 waigc=-2.737579e-012             paigc=-2.8389471e-019            aigsd=0.0049200857 laigsd=2.9842192e-011             waigsd=3.5714691e-011             paigsd=-2.7465182e-018 tvoff=0.000118118                ltvoff=1.92042e-010               wtvoff=1.43761e-010 ptvoff=-2.38008e-017              kt1=-0.21426871                lkt1=-4.7685822e-010 wkt1=3.6706608e-009             pkt1=-4.8542864e-016            kt2=-0.069985114 ute=-1.1281943                 lute=-3.2097168e-008            wute=-1.9818386e-008 pute=8.8588184e-015             ua1=1.5753978e-009             lua1=-1.2181818e-016 wua1=-8.3297292e-017            pua1=1.9066142e-023             ub1=-1.3720485e-018 lub1=1.5369671e-025             wub1=-4.856886e-026             pub1=1.0207212e-032 uc1=3.4801709e-010             luc1=-2.7125641e-017            wuc1=1.0801744e-017 puc1=1.4224686e-024             at=127861.76 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=4.3936792e-011             pcit=1.7827805e-017             lkt2=-6.6542211e-012 lat=-0.016924207               wat=-0.0016665178              pat=7.4493347e-010 wkt2=-4.1086466e-012            pkt2=1.836565e-018              u0_ff=4.97391e-05 u0_ss=8.01991e-05                u0_sf=4.97391e-05                u0_fs=8.01991e-05 lu0_ff=-2.63725e-11               lu0_ss=-2.26044e-11               lu0_sf=-2.63725e-11 lu0_fs=-2.26044e-11               wu0_ff=-3.00049e-11               wu0_ss=-7.09655e-12 wu0_sf=-3.00049e-11               wu0_fs=-7.09655e-12               pu0_ff=-3.95129e-18 pu0_ss=1.18539e-17                pu0_sf=-3.95129e-18               pu0_fs=1.18539e-17 vsat_mc=-2688.51                   lvsat_mc=0.000572652                wvsat_mc=0.000742028 pvsat_mc=-1.58052e-10               a0_ff=0.116903                   a0_ss=-0.22963 a0_sf=0.2                        a0_fs=-0.2                       la0_ff=3.46612e-08 la0_ss=-5.2e-13                   la0_sf=1.58e-13                   la0_fs=-1.58e-13 wa0_ff=3.79736e-08                wa0_ss=-1.94225e-08               wa0_sf=-5e-15 wa0_fs=5e-15                      pa0_ff=-3.95129e-15               pa0_ss=-1.4e-20 pa0_sf=7e-21                      pa0_fs=-7e-21                     at_mc=12098.3 lat_mc=-0.00257694                wat_mc=-0.00333913                pat_mc=7.11234e-10 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.25 pmos ( level=54                         lmin=9e-008                     lmax=2.16e-007 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.404469 lvth0=-1.1350568e-010            wvth0=-2.7229751e-010            pvth0=8.9879695e-017 k2=0.013420799                lk2=-4.1639477e-010            wk2=2.9456178e-009 pk2=-5.3514394e-017            cit=0.0024652488               wcit=5.6419786e-011 voff=-0.14471135                lvoff=-2.8442588e-009            wvoff=2.1019672e-009 pvoff=2.2789847e-016             eta0=0.13327531                 weta0=-9.0398552e-010 etab=-0.3320814                 wetab=8.7872798e-009             u0=0.015542008 lu0=1.6618663e-010             wu0=9.3033178e-011             pu0=-1.0959691e-017 ua=-4.0802569e-010            lua=-4.6504057e-017            wua=9.3851183e-018 pua=-2.4157659e-024            ub=1.1015376e-018             lub=-2.7280621e-026 wub=9.0855262e-026             pub=-5.2982959e-033            uc=1.8216748e-010 luc=-1.3959462e-017            wuc=-2.7465807e-018            puc=1.5739008e-025 vsat=57534.688                  lvsat=0.0040559479               wvsat=0.00098678605 pvsat=-3.2131678e-010            a0=-1.0276562                 la0=5.9972296e-008 wa0=6.0628344e-007             pa0=-9.559409e-014             ags=4.4897333 lags=-2.166068e-007             wags=-4.5388069e-007            pags=3.948762e-014 keta=0.052480379                lketa=-5.6935708e-009            wketa=2.3295106e-010 pketa=-1.8924007e-016            pclm=0.3879751                  lpclm=4.4357462e-009 wpclm=-1.6311615e-009            ppclm=-7.4040107e-016            pdiblc2=-0.00055555556 lpdiblc2=4.5755556e-010             wpdiblc2=7.907619e-010              ppdiblc2=-8.5693619e-017 aigbacc=0.014596901                laigbacc=-2.809567e-010             waigbacc=-4.2948696e-010 paigbacc=4.327135e-017              aigc=0.0059576279               laigc=-2.4487792e-012 waigc=-4.1876788e-012            paigc=2.4976548e-020             aigsd=0.0049660273 laigsd=2.0056632e-011             waigsd=3.2199665e-011             paigsd=-1.9978176e-018 tvoff=0.00104621                 ltvoff=-5.64211e-012              wtvoff=2.53501e-011 ptvoff=1.42066e-018               kt1=-0.2149209                 lkt1=-3.3794177e-010 wkt1=1.4313482e-009             pkt1=-8.4550466e-018            kt2=-0.070800257 ute=-1.3859295                 lute=2.2800429e-008             wute=3.2259386e-008 pute=-2.233747e-015             ua1=1.3047514e-009             lua1=-6.4170497e-017 wua1=2.0065461e-017             pua1=-2.9501244e-024            ub1=-9.1207945e-019 lub1=5.5723316e-026             wub1=-5.5910588e-026            pub1=1.1771e-032 uc1=2.729127e-010              luc1=-1.1128405e-017            wuc1=1.5066095e-017 puc1=5.1416171e-025             at=53080.956 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=-7.6097518e-011            pcit=-2.6847377e-018            lkt2=1.6697129e-010 lat=-0.00099589546             wat=0.0034889346               pat=-3.531779e-010 letab=1.2453137e-012             petab=-1.4196576e-019            leta0=5.29949e-010 peta0=-1.4626592e-016            wkt2=9.5707962e-011             pkt2=-1.9424373e-017 u0_ff=-0.000125221               u0_ss=-0.000109038               u0_sf=-0.000125221 u0_fs=-4.38267e-05               lu0_ff=1.08941e-11                lu0_ss=1.77031e-11 lu0_sf=1.08941e-11                lu0_fs=3.81298e-12                wu0_ff=-8.2082e-11 wu0_ss=6.19662e-11                wu0_sf=-8.2082e-11                wu0_fs=8.2082e-11 pu0_ff=7.14114e-18                pu0_ss=-2.85646e-18               pu0_sf=7.14114e-18 pu0_fs=-7.14114e-18               vsat_ff=1176.37                    vsat_ss=-1176.37 lvsat_ff=-0.000250566               lvsat_ss=0.000250566                wvsat_ff=-0.000134106 wvsat_ss=0.000134106                pvsat_ff=2.85645e-11                pvsat_ss=-2.85645e-11 a0_ff=0.403655                   a0_ss=-0.270546                  a0_sf=0.338095 a0_fs=-0.338095                  la0_ff=-2.64184e-08               la0_ss=8.71532e-09 la0_sf=-2.94143e-08               la0_fs=2.94143e-08                wa0_ff=3.2833e-08 wa0_ss=-4.62434e-08               wa0_sf=8e-15                      wa0_fs=-8e-15 pa0_ff=-2.85645e-15               pa0_ss=5.71291e-15                pa0_sf=2.1e-21 pa0_fs=-2.1e-21 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.26 pmos ( level=54                         lmin=5.4e-008                   lmax=9e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.39499874 lvth0=-9.3741874e-010            wvth0=2.0536969e-009             pvth0=-1.1248182e-016 k2=0.038029349                lk2=-2.5573386e-009            wk2=3.8528654e-010 pk2=1.6923442e-016             cit=-0.00031181049             wcit=2.5738886e-010 voff=-0.14976491                lvoff=-2.4045993e-009            wvoff=6.9174301e-009 pvoff=-1.9104681e-016            eta0=0.13054453                 weta0=-1.5029106e-010 etab=-0.67239289                wetab=1.5179788e-008             u0=0.017788866 lu0=-2.9290029e-011            wu0=-6.195608e-012             pu0=-2.3267867e-018 ua=-1.0769602e-009            lua=1.1693248e-017             wua=-3.970946e-017 pua=1.8554624e-024             ub=1.0635843e-018             lub=-2.3978677e-026 wub=6.0994231e-026             pub=-2.7003862e-033            uc=5.1677926e-011 luc=-2.6068709e-018            wuc=3.4595343e-018             puc=-3.8254193e-025 vsat=124385.32                  lvsat=-0.0017600574              wvsat=-0.0088172127 pvsat=5.3163111e-010             a0=11.450193                  la0=-1.0256006e-006 wa0=-1.4288424e-006            pa0=8.1461863e-014             ags=2 lags=0                          wags=0                          pags=0 keta=0.11931574                 lketa=-1.1508247e-008            wketa=-7.3319943e-009 pketa=4.6891018e-016             pclm=0.53023621                 lpclm=-7.9409705e-009 wpclm=-1.9117629e-008            ppclm=7.8092161e-016             pdiblc2=0.0042839506 lpdiblc2=3.6518519e-011             wpdiblc2=-4.6937037e-010            ppdiblc2=2.3937889e-017 aigbacc=0.0097606804               laigbacc=1.3979449e-010             waigbacc=3.17613e-010 paigbacc=-2.1726346e-017            aigc=0.0060755649               laigc=-1.2709297e-011 waigc=-4.5206742e-012            paigc=5.3947145e-020             aigsd=0.0051278845 laigsd=5.975051e-012              waigsd=8.7936375e-012             paigsd=3.8506727e-020 tvoff=-0.000198604               ltvoff=1.02657e-010               wtvoff=1.97805e-010 ptvoff=-1.3583e-017               kt1=-0.23099819                lkt1=1.0607826e-009 wkt1=1.3867019e-009             pkt1=-4.5708202e-018            kt2=-0.081462529 ute=-1.2708321                 lute=1.2786959e-008             wute=4.1362859e-008 pute=-3.0257492e-015            ua1=1.0810104e-009             lua1=-4.4705033e-017 wua1=-2.490834e-017             pua1=9.6259623e-025             ub1=-1.4142914e-018 lub1=9.9415756e-026             wub1=1.9460648e-025             pub1=-1.0023984e-032 uc1=5.9055556e-011             luc1=7.4771667e-018             wuc1=4.8215667e-017 puc1=-2.369851e-024             at=34172.706 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=1.6550664e-010             pcit=-2.0169047e-017            lkt2=1.094589e-009 lat=0.00064912223              wat=0.00039052345              pat=-8.361613e-011 letab=2.9608344e-008             petab=-5.562902e-016             leta0=7.675266e-010 peta0=-2.1183734e-016            wkt2=-3.0827166e-010            pkt2=1.5721855e-017 u0_ss=-0.000419753               u0_fs=-0.000498457               lu0_ss=4.47352e-11 lu0_fs=4.33657e-11                wu0_ss=2.49252e-10                wu0_fs=1.37574e-10 pu0_ss=-1.91503e-17               pu0_fs=-1.19689e-17               vsat_ff=-4117.28 vsat_ss=1703.7                     lvsat_ff=0.000209981                lvsat_ss=4.8e-10 wvsat_ff=0.00046937                 wvsat_ss=-0.000194222               pvsat_ff=-2.39379e-11 pvsat_ss=1.1e-17                    a0_ff=0.241666                   a0_ss=-0.411728 la0_ff=-1.2325e-08                la0_ss=2.09981e-08                wa0_ff=3.7e-14 wa0_ss=4.6937e-08                 pa0_ff=1.1e-21                    pa0_ss=-2.39379e-15 ua1_fs=-1.49537e-10               ua1_ss=-1.49537e-10               lua1_fs=1.30097e-17 lua1_ss=1.30097e-17                wua1_fs=4.12722e-17                wua1_ss=4.12722e-17 pua1_fs=-3.59068e-24               pua1_ss=-3.59068e-24 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.27 pmos ( level=54                         lmin=4.5e-008                   lmax=5.4e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.39627621 lvth0=-8.7226746e-010            wvth0=3.9160456e-009             pvth0=-2.074616e-016 k2=0.032122697                lk2=-2.2560993e-009            wk2=-1.5532523e-009 pk2=2.6809991e-016             cit=-0.0016586149              wcit=-5.0242539e-010 voff=-0.12711305                lvoff=-3.5598443e-009            wvoff=4.6691859e-009 pvoff=-7.6386352e-017            eta0=0.15960099                 weta0=-1.7298726e-009 etab=-0.38600244                wetab=2.0705904e-008             u0=0.022088483 lu0=-2.4857052e-010            wu0=-5.6845624e-010            pu0=2.6348506e-017 ua=-8.3669919e-010            lua=-5.6006523e-019            wua=-7.6229409e-017 pua=3.7179798e-024             ub=3.6683634e-019             lub=1.1555466e-026 wub=1.2799263e-025             pub=-6.1173045e-033            uc=-3.2490155e-011 luc=1.6857012e-018             wuc=1.9906236e-017             puc=-1.2213237e-024 vsat=31605.688                  lvsat=0.002971704                wvsat=0.0033508 pvsat=-8.8937537e-011            a0=-1.7883544                 la0=-3.5043467e-007 wa0=5.7840047e-007             pa0=-2.0907527e-014            ags=2 lags=0                          wags=0                          pags=0 keta=-0.41870493                lketa=1.5930807e-008             wketa=3.7472363e-008 pketa=-1.816112e-015             pclm=0.42637702                 lpclm=-2.6441516e-009 wpclm=-4.2778799e-009            ppclm=2.40944e-017               pdiblc2=0.00033333333 lpdiblc2=2.38e-010                  wpdiblc2=0                          ppdiblc2=0 aigbacc=0.018329406                laigbacc=-2.9721053e-010            waigbacc=-5.3316218e-010 paigbacc=2.1663188e-017             aigc=0.005980483                laigc=-7.8601224e-012 waigc=8.325656e-012              paigc=-6.012157e-019             aigsd=0.0049866545 laigsd=1.3177779e-011             waigsd=4.0425085e-011             paigsd=-1.5746971e-018 tvoff=0.00169607                 ltvoff=6.0287e-012                wtvoff=-1.49956e-010 ptvoff=4.15289e-018               kt1=-0.2588057                 lkt1=2.4789652e-009 wkt1=7.5334826e-009             pkt1=-3.1805664e-016            kt2=-0.06 ute=-0.64727531                lute=-1.9014437e-008            wute=-1.0180481e-007 pute=4.2758022e-015             ua1=1.8294851e-009             lua1=-8.287724e-017 wua1=-7.4435328e-017            pua1=3.4884726e-024             ub1=-1.2185786e-018 lub1=8.9434403e-026             wub1=6.0333651e-026             pub1=-3.1760703e-033 uc1=2.1811111e-010             luc1=-6.3466667e-019            wuc1=9.9053333e-018 puc1=-4.16024e-025              at=39857.423 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=2.3419366e-010             pcit=1.8581479e-017             lat=0.00035920165 wat=-0.0082634223              pat=3.577351e-010              letab=1.5002432e-008 petab=-8.3812212e-016            leta0=-7.1435259e-010            peta0=-1.3127868e-016 u0_fs=-0.000304943               u0_ss=0.000129015                lu0_fs=3.34963e-11 lu0_ss=1.6748e-11                 wu0_fs=8.41627e-11                wu0_ss=-3.56072e-11 pu0_fs=-9.24496e-18               pu0_ss=-4.62252e-18               vsat_ff=7950.62 vsat_ss=1703.7                     lvsat_ff=-0.000405481               lvsat_ss=4.8e-10 wvsat_ff=-0.00090637                wvsat_ss=-0.00019422                pvsat_ff=4.62249e-11 pvsat_ss=1.1e-17                    ua1_fs=2.69753e-10                ua1_ss=1.87654e-10 lua1_fs=-8.37412e-18               lua1_ss=-4.18702e-18               wua1_fs=-7.44519e-17 wua1_ss=-5.17929e-17               pua1_fs=2.31124e-24                pua1_ss=1.15562e-24 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model pch_lvt_mac.28 pmos ( level=54                         lmin=3.6e-08                    lmax=4.5e-008 wmin=1.08e-07                   wmax=2.7e-007                   vth0=-0.42924193 lvth0=5.1229258e-010             wvth0=8.2995035e-009             pvth0=-3.9156683e-016 k2=-0.0017061609              lk2=-8.3528729e-010            wk2=4.8310692e-010 pk2=1.8257282e-016             cit=-0.020938686               wcit=9.881098e-010 voff=-0.13912934                lvoff=-3.0551599e-009            wvoff=4.6540429e-010 pvoff=1.0017247e-016             eta0=0.15006173                 weta0=-1.1977037e-008 etab=-0.16299665                wetab=5.9608201e-009             u0=0.011691877 lu0=1.8808696e-010             wu0=3.673952e-010              pu0=-1.2957255e-017 ua=-1.1211106e-009            lua=1.1385215e-017             wua=4.7500881e-017 pua=-1.4786924e-024            ub=6.4165657e-019             lub=1.301661e-029 wub=-5.2285367e-026            pub=1.4543713e-033             uc=9.5351005e-011 luc=-3.6836275e-018            wuc=-2.6707209e-017            puc=7.3644097e-025 vsat=89657.737                  lvsat=0.00053351796              wvsat=0.00033937478 pvsat=3.7542324e-011             a0=12.6835                    la0=-9.5825256e-007 wa0=-1.4821903e-007            pa0=9.6104924e-015             ags=2 lags=0                          wags=0                          pags=0 keta=-0.20936152                lketa=7.1383838e-009             wketa=4.3595357e-008 pketa=-2.0732778e-015            pclm=-0.01580903                lpclm=1.5927662e-008 wpclm=7.3355932e-008             ppclm=-3.2365257e-015            pdiblc2=0.014827161 lpdiblc2=-3.7074074e-010            wpdiblc2=-1.4242963e-009            ppdiblc2=5.9820444e-017 aigbacc=0.01577298                 laigbacc=-1.8984062e-010            waigbacc=-7.3785619e-010 paigbacc=3.0260336e-017             aigc=0.0059246988               laigc=-5.5171827e-012 waigc=-8.7099292e-012            paigc=1.1427888e-019             aigsd=0.0057584583 laigsd=-1.9237981e-011            waigsd=-4.3425962e-011            paigsd=1.9470469e-018 tvoff=0.0071573                  ltvoff=-2.23343e-010              wtvoff=-6.68889e-010 ptvoff=2.59481e-017               kt1=0.12272755                 lkt1=-1.3545431e-008 wkt1=-3.9507918e-008            pkt1=1.6576822e-015             kt2=-0.10956788 ute=-1.5354099                 lute=1.8287215e-008             wute=4.9636726e-008 pute=-2.0847425e-015            ua1=1.2185202e-009             lua1=-5.7216715e-017 wua1=-1.0078675e-017            pua1=7.854932e-025              ub1=-3.1438447e-018 lub1=1.7029558e-025             wub1=2.8233965e-025             pub1=-1.2500322e-032 uc1=5.2688889e-010             luc1=-1.3603333e-017            wuc1=-2.5637333e-017 puc1=1.076768e-024              at=-37269.265 jtsswgs='7.8e-006*(1+0.3*iboffp_flag_lvt)'                                 jtsswgd='7.8e-006*(1+0.3*iboffp_flag_lvt)' lcit=1.0439567e-009             pcit=-4.4020998e-017            lkt2=2.081851e-009 lat=0.0035985226               wat=0.01163318                 pat=-4.7792219e-010 letab=5.6361885e-009             petab=-2.1882858e-016            leta0=-3.137037e-010 peta0=2.9910222e-016             wkt2=3.5607372e-009             pkt2=-1.4955096e-016 vth0_ss=-0.00516049                vth0_mc=0.0190123                  vth0_mcl=-0.0020642 lvth0_ss=2.16741e-10                lvth0_mc=-7.98516e-10               lvth0_mcl=8.66963e-11 wvth0_ss=1.4243e-09                 wvth0_mc=2.84859e-09                wvth0_mcl=5.69719e-10 pvth0_ss=-5.98204e-17               pvth0_mc=-1.19641e-16               pvth0_mcl=-2.39282e-17 cit_mcl=0.000387037                cit_mc=0.00774074                 wcit_mcl=-1.06822e-10 wcit_mc=-2.13644e-09               voff_mcl=-0.00937037                lvoff_mcl=3.93556e-10 wvoff_mcl=1.06822e-09                pvoff_mcl=-4.48653e-17               u0_ss=0.00272099 u0_fs=0.00100865                 u0_sf=-0.000774074               u0_mc=0.00258025 lu0_ss=-9.21148e-11               lu0_fs=-2.16741e-11               lu0_sf=3.25111e-11 lu0_mc=-1.0837e-10                wu0_ss=-7.50993e-10               wu0_fs=-2.78385e-10 wu0_sf=2.13644e-10                wu0_mc=-7.12148e-10               pu0_ss=2.54237e-17 pu0_fs=5.98206e-18                pu0_sf=-8.97307e-18               pu0_mc=2.99102e-17 vsat_fs=21864.2                    vsat_ff=-7950.62                   vsat_ss=7950.62 vsat_mc=8148.18                    vsat_mcl=-4237.01                   lvsat_fs=-0.000918296 lvsat_ff=0.00026237                 lvsat_ss=-0.00026237                lvsat_mc=-0.000342222 lvsat_mcl=0.000177956                wvsat_fs=-0.00249252                wvsat_ff=0.00090637 wvsat_ss=-0.00090637                wvsat_mc=-0.00427289                wvsat_mcl=-0.000854574 pvsat_fs=1.04686e-10                pvsat_ff=-2.99102e-11               pvsat_ss=2.99102e-11 pvsat_mc=1.79461e-10                pvsat_mcl=3.58923e-11                ua1_fs=3.28395e-10 ua1_ss=4.10494e-10                lua1_fs=-1.0837e-17                lua1_ss=-1.35463e-17 wua1_fs=-9.0637e-17                wua1_ss=-1.13296e-16               pua1_fs=2.99102e-24 pua1_ss=3.73878e-24                lcit_mcl=-1.62556e-11               lcit_mc=-3.25111e-10 pcit_mcl=4.48653e-18                pcit_mc=8.97307e-17 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_na_mac.global nmos ( modelid=13                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=1                          igbmod=1 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_na'              permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=1.96e-009                  toxm=1.96e-009                  dtox=3.3802e-010 epsrox=3.9                        toxref=3e-009                     wint=0 lint=0                          ll=0                          wl=0 lln=1                          wln=1                          lw=0 ww=0                          lwn=1                          wwn=1 lwl=0                          wwl=0                          llc=0 wlc=0                          lwc=0                          wwc=0 lwlc=0                          wwlc=0                          xl=-1.7e-008 xw=6e-009                     dlc=1.94e-008                  dwc=0 dlcig=2.5e-009                   xpart=1                          k1=0.033 k3=1                          k3b=-3.24                      w0=0 dvt0=0.13                       dvt1=0.1                        dvt2=0.1 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.56                       minv=-0.1                       voffl=0 dvtp0=2.5e-005                   dvtp1=0                          lpe0=2.3414e-006 lpeb=1e-007                     xj=6.7e-008                   ngate=2.106e+020 ndep=1e+016                     nsd=1e+020                     phin=0.15 cdsc=0                          cdscb=0                          cdscd=0 ud=0                          nfactor=1                          eta0=0.0030672 etab=0.2                        a1=0                          a2=1 b0=0                          b1=0                          dwg=0 dwb=0                          pdiblc1=0                          pdiblcb=1 drout=0.56                       pvag=0                          delta=0.01 pscbe1=1e+009                     pscbe2=1e-020                     fprout=500 pdits=0.065                      pditsd=0                          pditsl=0 rsh=18.0                       rdsw=120                        prwg=0 prwb=0                          wr=1                          alpha0=0 alpha1=4e-006                     beta0=2.4961                     agidl=1.85e-008 bgidl=2.3391e+009                cgidl=0.3                        egidl=0.27814 bigbacc=0.0005292                  cigbacc=0.82579                    nigbacc=3.7 aigbinv=0.2415                     bigbinv=0.0309                     cigbinv=0.006 eigbinv=1.1                        nigbinv=1                          bigc=0.0038588 cigc=0.21284                    bigsd=7.8302e-005                cigsd=2.1513e-020 nigc=7.9564                     poxedge=1                          pigcd=2.621 ntox=1                          vfbsdoff=0.01                       cgso=8.8e-011 cgdo=8.8e-011                   cgbo=0                          cgdl=3.0012e-010 cgsl=3.0012e-010                clc=0                          cle=0.6 cf='6.22e-011+9.73e-11*ccoflag_na'                                    ckappas=0.6 ckappad=0.6                        acde=0.29766                    moin=24 noff=4                          voffcv=-0.22327                   tvfbsdoff=0.01015 kt1l=0                          prt=0                          fnoimod=1 tnoimod=0                          em=1e+006                     ef=0.83 noia=0                          noib=0                          noic=0 lintnoi=-1.95e-009                 jss=2.76e-06                   jsd=2.76e-06 jsws=2.63e-12                   jswd=2.63e-12                   jswgs=2.63e-12 jswgd=2.63e-12                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=17.22                      bvd=17.22 xjbvs=1                          xjbvd=1                          jtsswgs=5.41e-008 jtsswgd=5.41e-008                  njtsswg=4.43                       xtsswgs=0.2348 xtsswgd=0.2348                     tnjtsswg=1                          vtsswgs=1.36 vtsswgd=1.36                       pbs=0.530                      pbd=0.530 cjs=0.000159                   cjd=0.000159                   mjs=0.336 mjd=0.336                      pbsws=0.4                        pbswd=0.4 cjsws=1.99e-010                  cjswd=1.99e-010                  mjsws=0.039 mjswd=0.039                      pbswgs=0.900                      pbswgd=0.900 cjswgs=1.49e-010                  cjswgd=1.49e-010                  mjswgs=0.500 mjswgd=0.500                      tpb=0.0023                     tcj=0.0022 tpbsw=0.0019                     tcjsw=0.00044                    tpbswg=0.004 tcjswg=0.003                      xtis=3                          xtid=3 dmcg=4.45e-008                  dmci=4.45e-008                  dmdg=0 dmcgt=0                          dwj=0                          xgw=0 xgl=2.64e-09                   rshg=16.42                      gbmin=1e-012 rbpb=50                         rbpd=50                         rbps=50 rbdb=50                         rbsb=50                         ngcon=1 xrcrg1=12                         xrcrg2=1 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.61 sigma_factor='sigma_factor_na' ccoflag='ccoflag_na' rcoflag='rcoflag_na' rgflag='rgflag_na' mismatchflag='mismatchflag_mos_na' globalflag='globalflag_mos_na' totalflag='totalflag_mos_na' global_factor='global_factor_na' local_factor='local_factor_na' sigma_factor_flicker='sigma_factor_flicker_na' noiseflag='noiseflagn_na' noiseflag_mc='noiseflagn_na_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w1='2.3875*0.35355' w2='0.70711*-0.35355' w3='0.54772*-0.0052117' w4='0.54772*-0.40307' w5='0.54772*-0.64548' w6='0.54772*-0.049915' w7='0.54772*-0.11513' w8='0.54772*-0.39385' w9='0' w10='0' tox_c='toxn_na'                  dxl_c='dxln_na'                  dxw_c='dxwn_na' cj_c='cjn_na'                   cjsw_c='cjswn_na'                 cjswg_c='cjswgn_na' cgo_c='cgon_na'                  cgl_c='cgln_na'                  ddlc_c='ddlcn_na' cf_c='cfn_na'                   dvth_c='dvthn_na'                 dlvth_c='dlvthn_na' dwvth_c='dwvthn_na'                dpvth_c='dpvthn_na'                du0_c='du0n_na' dlu0_c='dlu0n_na'                 dwu0_c='dwu0n_na'                 dpu0_c='dpu0n_na' dlk2_c='dlk2n_na'                 dwk2_c='dwk2n_na'                 dpk2_c='dpk2n_na' dvsat_c='dvsatn_na'                dlvsat_c='dlvsatn_na'               dwvsat_c='dwvsatn_na' dpvsat_c='dpvsatn_na'               dpdiblc2_c='dpdiblc2n_na'             dlpdiblc2_c='dlpdiblc2n_na' dwpdiblc2_c='dwpdiblc2n_na'            dppdiblc2_c='dppdiblc2n_na'            ntox_c='ntoxn_na' dags_c='dagsn_na'                 dlags_c='dlagsn_na'                dwags_c='dwagsn_na' dpags_c='dpagsn_na'                dua1_c='dua1n_na'                 monte_flag_c='monte_flagn_na' c1f_c='c1fn_na'                  c2f_c='c2fn_na'                  c3f_c='c3fn_na' global_mc='global_mc_flag_na' tox_g='toxn_na_ms_global'        dxl_g='dxln_na_ms_global'        dxw_g='dxwn_na_ms_global' cj_g='cjn_na_ms_global'         cjsw_g='cjswn_na_ms_global'       cjswg_g='cjswgn_na_ms_global' cgo_g='cgon_na_ms_global'        cgl_g='cgln_na_ms_global'        cf_g='cfn_na_ms_global' dvth_g='dvthn_na_ms_global'       dlvth_g='dlvthn_na_ms_global'      dwvth_g='dwvthn_na_ms_global' dpvth_g='dpvthn_na_ms_global'      du0_g='du0n_na_ms_global'        dlu0_g='dlu0n_na_ms_global' dwu0_g='dwu0n_na_ms_global'       dpu0_g='dpu0n_na_ms_global'       dvsat_g='dvsatn_na_ms_global' dwvsat_g='dwvsatn_na_ms_global'     dpdiblc2_g='dpdiblc2n_na_ms_global' ntox_g='ntoxn_na_ms_global'       dags_g='dagsn_na_ms_global'       dlags_g='dlagsn_na_ms_global' dwags_g='dwagsn_na_ms_global'      dua1_g='dua1n_na_ms_global' monte_flag_g='monte_flagn_na_ms_global'                                        ddlc_g='ddlcn_na_ms_global' weight1=-2.5235625 weight2=1.6628125 weight3=-0.642875 weight4=-0.625 weight5=-0.4297375 tox_1=8.388224e-012 tox_2=-1.2750464e-011 tox_3=-1.28768e-012 tox_4=4.797056e-011 tox_5=1.613696e-012 dxl_1=1.899264e-010 dxl_2=-2.886912e-010 dxl_3=-2.915456e-011 dxl_4=-1.0861184e-009 dxl_5=3.653632e-011 dxw_1=-8.181248e-010 dxw_2=-1.28768e-009 dxw_3=-2.892544e-010 dxw_4=-1.2013184e-024 dxw_5=-6.208512e-009 cj_1=1.3777e-006 cj_2=-5.38e-009 cj_3=2.7027e-008 cj_4=-1.5241e-022 cj_5=-1.7865e-007 cjsw_1=1.7242e-012 cjsw_2=-6.7335e-015 cjsw_3=3.3826e-014 cjsw_4=9.728e-028 cjsw_5=-2.236e-013 cjswg_1=1.291e-012 cjswg_2=-5.0416e-015 cjswg_3=2.5327e-014 cjswg_4=3.4927e-028 cjswg_5=-1.6742e-013 cgo_1=-7.6248e-013 cgo_2=2.9776e-015 cgo_3=-1.4958e-014 cgo_4=-4.0643e-028 cgo_5=9.8877e-014 cgl_1=-2.6004e-012 cgl_2=1.0155e-014 cgl_3=-5.1015e-014 cgl_4=-1.3907e-027 cgl_5=3.3722e-013 cf_1=-5.3894e-013 cf_2=2.1046e-015 cf_3=-1.0573e-014 cf_4=-1.5443e-028 cf_5=6.9888e-014 dvth_1=0.00650496 dvth_2=0.00418845 dvth_3=0.00091119 dvth_4=-2.53428e-018 dvth_5=-0.001777965 dlvth_1=4.118345e-010 dlvth_2=2.85247e-010 dlvth_3=-1.320215e-012 dlvth_4=1.022105e-025 dlvth_5=-1.124135e-010 dwvth_1=3.0902e-010 dwvth_2=-7.9675e-010 dwvth_3=-1.6281e-010 dwvth_4=7.2642e-025 dwvth_5=1.3248e-010 dpvth_1=4.9554e-020 dpvth_2=1.7632e-016 dpvth_3=6.648e-017 dpvth_4=-2.8372e-031 dpvth_5=-3.9575e-017 du0_1=0.00057603 du0_2=0.00098093 du0_3=0.00021155 du0_4=-3.2076e-019 du0_5=-0.00028695 dlu0_1=1.2431e-011 dlu0_2=1.228e-010 dlu0_3=3.4787e-011 dlu0_4=-1.6778e-025 dlu0_5=-2.8644e-011 dwu0_1=5.821e-011 dwu0_2=-2.176e-011 dwu0_3=-3.195e-011 dwu0_4=1.2893e-025 dwu0_5=-1.5767e-012 dpu0_1=-1.8369e-017 dpu0_2=3.9488e-017 dpu0_3=1.5769e-017 dpu0_4=-5.9128e-032 dpu0_5=-6.5395e-018 dvsat_1=15.77 dvsat_2=7508.8 dvsat_3=-5708.3 dvsat_4=2.0945e-011 dvsat_5=-1297.4 dvsat_max=-28000 dwvsat_1=-1.5325e-006 dwvsat_2=-0.00012237 dwvsat_3=0.00089041 dwvsat_4=-3.2029e-018 dwvsat_5=-1.5081e-005 dpdiblc2_1=-0.00024756 dpdiblc2_2=9.6676e-007 dpdiblc2_3=-4.8566e-006 dpdiblc2_4=-9.8936e-020 dpdiblc2_5=3.2103e-005 ntox_1=-0.066244 ntox_2=0.00014425 ntox_3=0.0066772 ntox_4=-9.6357e-018 ntox_5=0.0075346 dags_1=0.01426 dags_2=-8.4785e-005 dags_3=0.0023077 dags_4=-1.5633e-017 dags_5=-0.0021177 dlags_1=-1.2378e-008 dlags_2=4.8338e-011 dlags_3=-2.4283e-010 dlags_4=3.3413e-023 dlags_5=1.6052e-009 dwags_1=-1.8653e-009 dwags_2=1.6983e-011 dwags_3=-7.1259e-010 dwags_4=2.4825e-024 dwags_5=3.3136e-010 dua1_1=2.4756e-011 dua1_2=-9.6676e-014 dua1_3=4.8566e-013 dua1_4=-5.2172e-027 dua1_5=-3.2103e-012 monte_flag_1=0.12365 monte_flag_2=-0.18795 monte_flag_3=-0.0189808 monte_flag_4=-0.707108 monte_flag_5=0.0237867 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.994 b_4=0.001185                   c_4=-0.04648                   d_4=0.007355 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0.000005                   g_4_2=-1.8555e-08 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.00662                    mis_a_2=0.55                       mis_a_3=0.04146 mis_b_1=0.0035                     mis_b_2=0                          mis_b_3=-0.1 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.0007                     mis_d_2=0                          mis_d_3=0 mis_e_1=0.025                      mis_e_2=0.6                        mis_e_3=0.06 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-1.7e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0                       bidirectionflag=1 designflag=1 cf0=6.22e-011                  cco=9.73e-11 noimod=1                          noic2='2.236'                    noic3='0.6' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.453e-6            sbref0=0.453e-6 samax=10e-6		sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=1                   lreflod=0.9e-6              llodref=2 lod_clamp=-1e90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=0 kvth00=-0e-9               lkvth00=0e-8                wkvth00=0e-8 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0e-11 lodeta00=1 wlod00=0 ku000=-0e-9               lku000=0e-28               wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0.0e-8              lkvth000=0e-23               wkvth000=-0e-16         	pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=0.27e-6 ku01=-1e-7               lku01=0.8e-13                   wku01=3e-14 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=-3.5 kvth01=10e-8                lkvth01=-40e-15            wkvth01=-1.0e-14 pkvth01=0                   llodvth1=1                   wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.0              lku02=0e-8              wku02=0e-8 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=-4 kvth02=5e-2              lkvth02=5.5e-7               wkvth02=-5e-8 pkvth02=0.0e-15             llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0 lodeta02=1 wlod02=0 ku002=-0.1                   lku002=-0e-10              wku002=0e-9         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0e-3                lkvth002=0e-18               wkvth002=0e-9         	    pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=-0.04              lku03=-0.6e-8             wku03=10e-8 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=-3.4 kvth03=15.0e-3              lkvth03=1e-9                wkvth03=5.0e-10 pkvth03=0e-16               llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=0                   lku003=-1.3e-8                   wku003=2e-9         		pku003=10e-16 llodku003=1                   wlodku003=1 kvth003=0e-3                lkvth003=-0e-9               wkvth003=0e-10         	pkvth003=-0e-18 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=1.e-7             sa_b1=0.99e-7             dpdbinflag=1 w_b=9e-6                w_b1=10e-6 sparef=1.54e-7             spamax=4.8e-7              spamin=1.54e-7 kvth0dpc='10.4'                 wkvth0dpc='-1.8e-6'              wdpckvth0=1 lkvth0dpc='1.2e-8'              ldpckvth0=1                   pkvth0dpc='10e-15*0' ku0dpc='-1.0'                 wku0dpc='2.8e-7*1'           wdpcku0=1 lku0dpc='0.2e-7'            ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc='2.5*0'               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc='2'                wdpc=0 kvth0dpc_b1=-0.0            kvth0dpc_b2=-0.0          dpcbinflg=1 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0  kvth0dpl='-30.0'                   wkvth0dpl='4e-7*0+5e-6'            wdplkvth0=1  lkvth0dpl='-0e-7'         ldplkvth0='1.0'               pkvth0dpl=0.00e+00  ku0dpl='2'                  wku0dpl='7e-7*0'             wdplku0=1  lku0dpl='-2e-7'              ldplku0='1.0'                 pku0dpl='2e-13*0'  keta0dpl='0'                 wketa0dpl=0.00e+00            wdplketa0=1  kvsatdpl=1                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000           dplbinflg=1 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx='-0.1*0'              wkvth0dpx='1e-6*0'               wdpxkvth0=1 lkvth0dpx='1e-7*0'              ldpxkvth0=1.0                 pkvth0dpx='8e-14*0' ku0dpx='-0.4'                wku0dpx=1e-6                wdpxku0=1 lku0dpx=0e-8              ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=-3                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000          dpxbinflg=1 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0                wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps=-0                 wku0dps=-0.0e-9             wdpsku0=1 lku0dps=0.0e-16             ldpsku0=1.0                 pku0dps=0.0e-23 keta0dps=0.00                wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000           dpsbinflg=1 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0  kvth0dpa='-0.12'             wkvth0dpa='-0e-08'            wdpakvth0=1  lkvth0dpa=0.00e+00           ldpakvth0=1                   pkvth0dpa=0.00e+00  ku0dpa=-0.0                     wku0dpa=0.0e-9              wdpaku0=1  lku0dpa='-0.0e-08'           ldpaku0=1                     pku0dpa=0.00e+00  keta0dpa=0                   wketa0dpa=0.00e+00            wdpaketa0=1  ka0dpa=0                     wka0dpa=0                     wdpaka0=1  lka0dpa=0.00e+00             ldpaka0=1                     pka0dpa=0.00e+00  kvsatdpa=0                   wdpa=0 kvth0dpa_b1=0.000             kvth0dpa_b2='-0.02'           dpabinflg=1 ku0dpa_b1=-0.00             ku0dpa_b2='0.05*0' keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.08e-7             spbmax='4.8e-7+6.8e-7'     spbmin='1.54e-7+3.54e-7' pse_mode=1 kvth0dp2=0              	 wkvth0dp2=0            		 wdp2kvth0=1 lkvth0dp2=0e-8           	 ldp2kvth0=1                   pkvth0dp2=0 ku0dp2=0             	     wku0dp2=0e-9             	 wdp2ku0=1 lku0dp2=0.0e-8          	 ldp2ku0=1                 	 pku0dp2=0 keta0dp2=0               	 wketa0dp2=0               	 wdp2keta0=1 kvsatdp2=0.0               	 wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0                kvth0dp2l_b2=0                dp2lbinflg=0 ku0dp2l_b1=0                ku0dp2l_b2=0 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=1.0                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1e-7 kvth0enx=-0.02            	 wkvth0enx=-1.2e-5             wenxkvth0=0.5 lkvth0enx=0          		 lenxkvth0=1                   pkvth0enx=-0.3e-12 ku0enx=-2.5         		 wku0enx=-2.5e-4      		 wenxku0=0.5 lku0enx=10e-8          	 lenxku0=1                   pku0enx=-5e-12 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0                   wka0enx=0                   wenxka0=1 lka0enx=0          		 lenxka0=1                   pka0enx=0 kvsatenx=0.6                 wenx=0                   ku0enx0=0 eny0=2e-6 enyref=2e-6             enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0.007          	 wkvth0eny=0       		     wenykvth0=1 lkvth0eny=0        			 lenykvth0=1                   pkvth0eny=2.5e-17 ku0eny=20          		 wku0eny=2e-8        		 wenyku0=1 ku0eny0=0.00          		 wku0eny0=0                   weny0ku0=1 lku0eny=8e-6       		 lenyku0=1                 	 pku0eny=2e-16 keta0eny=0               	 wketa0eny=0                   wenyketa0=1 ka0eny=0              	 wka0eny=0             		 wenyka0=1 lka0eny=0      		     lenyka0=1                	 pka0eny=0 kvsateny=0.5               	 weny=0 kvth0eny1=-4.5e-4          	 wkvth0eny1=0        		     weny1kvth0=1 lkvth0eny1=0             	 leny1kvth0=1                  pkvth0eny1=-1e-18 ku0eny1=-0.005        	 wku0eny1=-0e-9            	 weny1ku0=1 lku0eny1=0e-4      		 leny1ku0=0.5                pku0eny1=-0.4e-12 keta0eny1=0              	 wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1                	 pka0eny1=0 kvsateny1=0.5                weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.8126e-5           ringxmin=0 kvth0rx=0.00              	 wkvth0rx=0e-9          	     wrxkvth0=1 lkvth0rx=0              	 lrxkvth0=1                	 pkvth0rx=0e-16 ku0rx=1.2              	 wku0rx=10e-8           	 wrxku0=1 lku0rx=0e-9        		 lrxku0=1                   pku0rx=0 keta0rx=0                	 wketa0rx=0                   wrxketa0=1 kvsatrx=0.1                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=1.6027e-5           ringymin=0 kvth0ry=-0.005           	 wkvth0ry=0           	     wrykvth0=1 lkvth0ry=0              	 lrykvth0=1                 	 pkvth0ry=0 ku0ry=-0.15          	 wku0ry=0           		 wryku0=1 lku0ry=0        			 lryku0=1                 	 pku0ry=0 keta0ry=0                	 wketa0ry=0                   wryketa0=1 kvsatry=0.5                 wry=0 kvth0ry0=0                	 ku0ry0=0 sfxref=8.26e-7           sfxmax=10e-6              minwodx=0.0e-6 sfxmin=0.252e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-2.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=0.00              lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0009           lkvth0odx1b=-0.2e-9            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.007            lku0odx1b=0                 lodx1bku0=1.0 wku0odx1b=-0.0e-5           wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6 sfymax=10e-6             minwody=0.9e-6            wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-1.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.000            lkvth0odyb=0.0e-10           lodybkvth0=1.0 wkvth0odyb=-2.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=-0.03             lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-1.0e-7           wodybku0=1.0               pku0odyb=0 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=0 oseflag=1 wpeflag=0 )
.model nch_na_mac.1 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=9e-007                     wmax=9.01e-06                   vth0=-0.0068103451 lvth0=-3.5260427e-009            wvth0=-3.5323123e-009            pvth0=1.0222853e-015 k2=0.0028049942               lk2=-1.9512986e-009            wk2=-4.0032633e-009 pk2=6.7091617e-016             cit=0.0013297044               lcit=1.033371e-009 wcit=-4.4686001e-010            pcit=3.9457739e-016             voff=-0.14766073 lvoff=-1.4218989e-08             wvoff=-1.1778021e-09             pvoff=-2.9776381e-15 u0=0.057589269                lu0=4.3988685e-009             wu0=-2.006473e-009 pu0=1.7717156e-015             ua=-9.6255495e-011            lua=1.3285659e-016 wua=-7.4330584e-018            pua=-6.5730711e-023            ub=3.7193439e-018 lub=-5.9569107e-025            wub=-1.4112208e-025            pub=2.1350104e-031 uc=-1.0073287e-011            luc=6.5834094e-019             wuc=6.6002655e-019 puc=-5.9290185e-024            vsat=87310.325                  lvsat=0.067038848 wvsat=-0.00220844                pvsat=2.1684395e-008             a0=12.183784 la0=-6.442046e-006             wa0=3.4403788e-006             pa0=-2.1483752e-012 ags=1.4905331                  lags=5.5944125e-006             wags=-1.9898461e-007 pags=-1.6060373e-012            keta=-0.037215497               lketa=-3.6877987e-008 wketa=2.3285769e-009             pketa=-1.0168102e-014            pclm=1.2745396 lpclm=2.2871112e-007             wpclm=3.2943676e-008             ppclm=-2.9593304e-013 pdiblc2=0.015257958                lpdiblc2=1.5146383e-008             wpdiblc2=-4.8722199e-010 ppdiblc2=8.9011727e-015             aigbacc=0.020554714                laigbacc=-9.3156101e-009 waigbacc=-8.0252361e-009            paigbacc=8.0424737e-015             aigc=0.011541324 laigc=-1.9968149e-010            waigc=1.0383346e-011             paigc=-1.4576083e-017 aigsd=0.0085202601               laigsd=3.5530611e-010             waigsd=4.1885437e-012 paigsd=-7.2237256e-020            tvoff=0.00423599                 ltvoff=-2.88498e-010 wtvoff=-6.68345e-011              ptvoff=-5.69723e-016              kt1=-0.27150765 lkt1=5.3613682e-009             wkt1=-1.5400935e-008            pkt1=3.8501639e-015 kt2=-0.014492425               lkt2=5.1507882e-010             wkt2=-2.2074476e-009 pkt2=1.876454e-015              ute=-2.0129581                 lute=1.0147027e-006 wute=-2.503939e-008             pute=2.2492884e-013             ua1=2.7647275e-009 lua1=2.1619422e-015             wua1=2.1058001e-016             pua1=3.9124865e-022 ub1=-5.8946861e-018            lub1=1.5180406e-024             wub1=-5.446458e-025 pub1=7.3532224e-031             uc1=6.5483307e-011             luc1=1.8827938e-017 wuc1=-3.5748801e-017            puc1=3.1566191e-023             at=101216.32 pat=9.8620157e-08              wat=-0.010966325               lat=-0.010938349 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na_mac.2 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=-0.026553619 lvth0=1.3907268e-008             wvth0=-1.2644318e-009            pvth0=-9.8025314e-016 k2=0.0010363134               lk2=-3.895534e-010             wk2=-3.6523877e-009 pk2=3.6109295e-016             cit=0.0023075556               lcit=1.6992844e-010 voff=-0.13609383                lvoff=-2.4432557e-008            wvoff=-1.3959858e-008 pvoff=8.308917e-015              u0=0.05871041                 lu0=3.4089013e-009 wu0=7.938624e-011              pu0=-7.009801e-017             ua=2.2792048e-010 lua=-1.5339079e-016            wua=-7.791867e-017             pua=-3.4919154e-024 ub=3.0494108e-018             lub=-4.1401444e-027            wub=5.8441792e-026 pub=3.728614e-032              uc=-5.0326428e-012            luc=-3.7925483e-018 wuc=-1.5185732e-017            puc=8.0627865e-024             vsat=129558.38 lvsat=0.029733819                wvsat=0.051026787                pvsat=-2.5322311e-008 a0=3.8182996                  la0=9.4467628e-007             wa0=1.9766206e-006 pa0=-8.5587671e-013            ags=6.6401707                  lags=1.0472825e-006 wags=-3.5015507e-006            pags=1.3101286e-012             keta=-0.10274653 lketa=2.0985916e-008             wketa=-5.6689725e-010            pketa=-7.6113978e-015 pclm=1.6345456                  lpclm=-8.9174231e-008            wpclm=-3.4514056e-007 ppclm=3.7915338e-014             pdiblc2=0.028318788                lpdiblc2=3.613669e-009 wpdiblc2=1.5916498e-008             ppdiblc2=-5.5833117e-015            aigbacc=0.010338038 laigbacc=-2.9428497e-010            waigbacc=1.1889276e-009             paigbacc=-9.3632912e-017 aigc=0.011446371                laigc=-1.1583827e-010            waigc=-2.0789262e-011 paigc=1.2949329e-017             aigsd=0.008775799                laigsd=1.2966528e-010 waigsd=4.0912263e-012             paigsd=1.3694027e-020             tvoff=0.00490227 ltvoff=-8.76821e-010              wtvoff=-9.2206e-010               ptvoff=1.85441e-016 kt1=-0.24562571                lkt1=-1.749238e-008             wkt1=-1.1887319e-008 pkt1=7.4764083e-016             kt2=-0.013213976               lkt2=-6.1379164e-010 wkt2=1.2737189e-010             pkt2=-1.8519161e-016            ute=-0.87350136 lute=8.562367e-009              wute=5.6824425e-007             pute=-2.9894062e-013 ua1=5.6262219e-009             lua1=-3.6475736e-016            wua1=2.400698e-015 pua1=-1.5426256e-021            ub1=-4.5452813e-018            lub1=3.2651617e-025 wub1=-8.4807482e-025            pub1=1.0032501e-030             uc1=9.0378549e-011 luc1=-3.1545605e-018            wuc1=-3.2174373e-017            puc1=2.8409971e-023 at=183856.3                   lat=-0.08390946                wat=0.14796664 pat=-4.1717652e-08 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na_mac.3 nmos ( level=54                         lmin=2.7e-07                    lmax=4.5e-007 wmin=9e-007                     wmax=9.01e-06                   vth0=0.012084072 lvth0=-2.822852e-009             wvth0=-2.5212515e-008            pvth0=9.3892669e-015 k2=0.00060357882              lk2=-2.0217934e-010            wk2=-2.9806109e-009 pk2=7.0213607e-017             cit=0.0022783333               lcit=1.8258167e-010 voff=-0.17537502                lvoff=-7.4238045e-009            wvoff=2.2065957e-008 pvoff=-7.2902609e-015            u0=0.074560156                lu0=-3.4540388e-009 wu0=-3.400348e-010             pu0=1.115113e-016              ua=2.4388379e-010 lua=-1.6030291e-016            wua=-1.9019735e-017            pua=-2.8995155e-023 ub=3.3917291e-018             lub=-1.5236395e-025            wub=3.477302e-025 pub=-8.7975741e-032            uc=1.3059475e-011             luc=-1.1626435e-017 wuc=-3.0638179e-018            puc=2.8139976e-024             vsat=195736.64 lvsat=0.0010786294               wvsat=-0.017931732               pvsat=4.5367281e-009 a0=13.027778                  la0=-3.0430278e-006            ags=12.267075 lags=-1.3891669e-006            wags=-3.9764208e-006            pags=1.5157474e-012 keta=-0.1104894                 lketa=2.4338578e-008             wketa=-4.0889516e-008 pketa=9.8482962e-015             pclm=2.3121335                  lpclm=-3.8256977e-007 wpclm=-6.1961403e-007            ppclm=1.5676235e-013             pdiblc2=0.030246782 lpdiblc2=2.7788479e-009             wpdiblc2=2.2844182e-008             ppdiblc2=-8.5829991e-015 aigbacc=0.00950659                 laigbacc=6.5731925e-011             waigbacc=2.3398487e-009 paigbacc=-5.9198171e-016            aigc=0.011258525                laigc=-3.4501068e-011 waigc=6.7787173e-011             paigc=-2.5404267e-017            aigsd=0.0090752601 laigsd=-1.3903391e-015            waigsd=4.152543e-012              paigsd=-1.2856107e-020 tvoff=0.0037668                  ltvoff=-3.85164e-010              wtvoff=-5.28698e-010 ptvoff=1.51154e-017               kt1=-0.26685297                lkt1=-8.3009782e-009 wkt1=-3.1131592e-008            pkt1=9.0804109e-015             kt2=-0.013965575 lkt2=-2.8834928e-010            wkt2=-9.7863456e-010            pkt2=2.9370919e-016 ute=-1.1347351                 lute=1.2167659e-007             wute=-2.9383808e-007 pute=7.4341034e-014             ua1=5.3402563e-009             lua1=-2.4093427e-016 wua1=-2.4887582e-015            pua1=5.7450896e-022             ub1=-5.2989451e-018 lub1=6.5285262e-025             wub1=3.5335204e-024             pub1=-8.9398067e-031 uc1=1.3474436e-010             luc1=-2.2364958e-017            wuc1=5.9490272e-017 puc1=-1.128082e-023             at=70412.693                  lat=-0.034788374 wat=0.072394591                pat=-8.9949544e-009 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na_mac.4 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.016899424 lvth0=2.0636588e-009             wvth0=5.6083935e-009             pvth0=-4.0419843e-015 k2=0.0016772161               lk2=-3.0471121e-009            wk2=-2.9814964e-009 pk2=1.6637232e-015             cit=0.00083648148              lcit=1.4688869e-009 voff=-0.13896204                lvoff=-3.9331792e-008            wvoff=-9.0588147e-009 pvoff=1.9774561e-014             u0=0.055374619                lu0=6.3544045e-009 ua=-6.9385657e-011            lua=1.58746e-018               wua=-3.1777132e-017 pua=5.3199121e-023             ub=3.5469249e-018             lub=-2.1042608e-025 wub=1.5089507e-026             pub=-1.3554904e-031            uc=-7.3590206e-012 luc=-2.3723918e-017            wuc=-1.7990992e-018            puc=1.6161308e-023 vsat=83566.603                  lvsat=0.1027062                  wvsat=0.0011833715 pvsat=-1.0630226e-008            a0=16.734574                  la0=-1.1085689e-005 wa0=-6.8263761e-007            pa0=2.0587654e-012             ags=1.1105954 lags=5.3737893e-006             wags=1.4523889e-007             pags=-1.4061526e-012 keta=-0.019875054               lketa=-5.6231503e-008            wketa=-1.3381864e-008 pketa=7.3661845e-015             pclm=1.3411741                  lpclm=-3.6986734e-007 wpclm=-2.7427256e-008            ppclm=2.4637904e-013             pdiblc2=-0.00013013477 lpdiblc2=1.5317226e-008             wpdiblc2=1.345439e-008              ppdiblc2=8.7463888e-015 aigbacc=0.012571479                laigbacc=-1.2110156e-009            waigbacc=-7.9242481e-010 paigbacc=6.9971111e-016             aigc=0.011572639                laigc=-2.4646096e-010 waigc=-1.7988186e-011            paigc=2.7806116e-017             aigsd=0.0085204535 laigsd=3.5510596e-010             waigsd=4.0133219e-012             paigsd=1.0910111e-019 tvoff=0.00466965                 ltvoff=-1.21379e-009              wtvoff=-4.5973e-010 ptvoff=2.68595e-016               kt1=-0.28366974                lkt1=2.4027924e-008 wkt1=-4.3820765e-009            pkt1=-1.3061736e-014            kt2=-0.019689067 lkt2=5.0234461e-009             wkt2=2.5007098e-009             pkt2=-2.2081268e-015 ute=-2.0356833                 lute=1.218843e-006              wute=-4.4503757e-009 pute=3.9977725e-014             ua1=2.6080232e-009             lua1=4.4210113e-015 wua1=3.5255411e-016             pua1=-1.655468e-021             ub1=-5.6895078e-018 lub1=-1.6465438e-024            wub1=-7.3053731e-025            pub1=3.6024357e-030 uc1=7.8724263e-011             luc1=1.6250883e-017             wuc1=-4.7745107e-017 puc1=3.3901003e-023             at=80855.631                  pat=-6.7271761e-08 wat=0.0074804579               lat=0.17216531                 wu0=0 pu0=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na_mac.5 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.034601982 lvth0=1.7695017e-008             wvth0=6.0273849e-009             pvth0=-4.4119537e-015 k2=-0.0023620572              lk2=5.1956623e-010             wk2=-5.7346397e-010 pk2=-4.6256943e-016            cit=0.0023075556               lcit=1.6992844e-010 voff=-0.16512833                lvoff=-1.6226959e-008            wvoff=1.2345394e-008 pvoff=8.7464518e-016             u0=0.057923726                lu0=4.1035426e-009 wu0=7.921211e-010              pu0=-6.99443e-016              ua=7.8976859e-011 lua=-1.2941664e-016            wua=5.7024248e-017             pua=-2.5212497e-023 ub=3.15788e-018               lub=1.3310059e-025             wub=-3.9831304e-026 pub=-8.7053969e-032            uc=-6.045637e-011             luc=2.3161042e-017 wuc=3.5028165e-017             puc=-1.6357166e-023            vsat=194796.32 lvsat=0.0044903591               wvsat=-0.0080787919              pvsat=-2.4517361e-009 a0=0.050857474                la0=3.6460328e-006             wa0=5.3899231e-006 pa0=-3.3033058e-012            ags=4.6383254                  lags=2.2588037e-006 wags=-1.6878789e-006            pags=2.1249041e-013             keta=-0.10603412 lketa=1.9846953e-008             wketa=2.4116593e-009             pketa=-6.5794968e-015 pclm=1.2277814                  lpclm=-2.6974158e-007            wpclm=2.3387793e-008 ppclm=2.0150936e-013             pdiblc2=0.021241642                lpdiblc2=-3.5540534e-009 wpdiblc2=2.2328392e-008             ppdiblc2=9.1064483e-016             aigbacc=0.012333305 laigbacc=-1.0007086e-009            waigbacc=-6.1878471e-010            paigbacc=5.463869e-016 aigc=0.011405696                laigc=-9.9050123e-011            waigc=1.6062607e-011 paigc=-2.2607342e-018            aigsd=0.008775738                laigsd=1.2968976e-010 waigsd=4.1464915e-012             paigsd=-8.4876769e-021            tvoff=0.00499287 ltvoff=-1.4992e-009               wtvoff=-1.00415e-009              ptvoff=7.49315e-016 kt1=-0.21240461                lkt1=-3.8899183e-008            wkt1=-4.1985633e-008 pkt1=2.0142204e-014             kt2=-0.014003022               lkt2=2.6683651e-012 wkt2=8.4224731e-010             pkt2=-7.4370437e-016            ute=0.26067566 lute=-8.0884198e-007            wute=-4.5932013e-007            pute=4.4162772e-013 ua1=1.2578332e-008             lua1=-4.3827714e-015            wua1=-3.8979137e-015 pua1=2.0976952e-021             ub1=-1.1883012e-017            lub1=3.8223209e-024 wub1=5.7999097e-024             pub1=-2.163949e-030             uc1=2.6678564e-011 luc1=6.2207235e-017             wuc1=2.5537813e-017             puc1=-3.0807815e-023 at=508696.69                  lat=-0.20561834                wat=-0.14633874 pat=6.8550591e-08 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na_mac.6 nmos ( level=54                         lmin=2.7e-07                    lmax=4.5e-007 wmin=5.4e-007                   wmax=9e-007                     vth0=-0.040881325 lvth0=2.0413973e-008             wvth0=2.2774135e-008             pvth0=-1.1663296e-014 k2=0.0017556588               lk2=-1.2634048e-009            wk2=-4.0243954e-009 pk2=1.0316839e-015             cit=0.0054759722               lcit=-1.201996e-009 wcit=-2.8970608e-009            pcit=1.2544273e-015             voff=-0.17090462 lvoff=-1.3725825e-08             wvoff=1.8015776e-08              pvoff=-1.5806303e-15 u0=0.076583782                lu0=-3.9762615e-009            wu0=-2.1734402e-009 pu0=5.846451e-016              ua=3.84221e-010               lua=-2.6158736e-016 wua=-1.4616525e-016            pua=6.2768557e-023             ub=4.039064e-018 lub=-2.4845206e-025            wub=-2.3875522e-025            pub=-9.1991338e-034 uc=2.5501667e-011             luc=-1.4058788e-017            wuc=-1.4336443e-017 puc=5.0177094e-024             vsat=195118.82                  lvsat=0.0043507182 wvsat=-0.017371983               pvsat=1.5722156e-009             a0=26.234148 la0=-7.6913318e-006            wa0=-1.1964971e-005            pa0=4.2113635e-012 ags=6.7931405                  lags=1.3257688e-006             wags=9.8296353e-007 pags=-9.4398437e-013            keta=-0.18203503                lketa=5.2755346e-008 wketa=2.3930824e-008             pketa=-1.5897295e-014            pclm=0.33048768 lpclm=1.1878662e-007             wpclm=1.1757571e-006             ppclm=-2.9746654e-013 pdiblc2=0.005514413                lpdiblc2=3.2558369e-009             wpdiblc2=4.5251708e-008 ppdiblc2=-9.0151512e-015            aigbacc=0.011289018                laigbacc=-5.4853213e-010 waigbacc=7.2496905e-010             paigbacc=-3.545848e-017             aigc=0.011346511 laigc=-7.3423325e-011            waigc=-1.1928228e-011            paigc=9.8592971e-018 aigsd=0.0090753192               laigsd=-2.8890709e-014            waigsd=4.0990391e-012 paigsd=1.2059228e-020             tvoff=0.00254742                 ltvoff=-4.40321e-010 wtvoff=5.76053e-010               ptvoff=6.50882e-017               kt1=-0.37467001 lkt1=3.1361735e-008             wkt1=6.6550652e-008             pkt1=-2.6854007e-014 kt2=-0.012926071               lkt2=-4.6365121e-010            wkt2=-1.920425e-009 pkt2=4.5253274e-016             ute=-3.4173416                 lute=7.8373951e-007 wute=1.7742034e-006             pute=-5.2548798e-013            ua1=1.4081773e-009 lua1=4.5390557e-016             wua1=1.0737054e-015             pua1=-5.5015938e-023 ub1=-8.285083e-018             lub1=2.2644174e-024             wub1=6.2389614e-024 pub1=-2.3540583e-030            uc1=2.3881436e-010             luc1=-2.9647565e-017 wuc1=-3.4797147e-017            puc1=-4.6827773e-024            at=157086.28 lat=-0.053371032               wat=-0.00613168                pat=7.840933e-09 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na_mac.7 nmos ( level=54                         lmin=9e-007                     lmax=9.01e-06 wmin=4.5e-07                    wmax=5.4e-007                   vth0=-0.03684026 lvth0=2.0512991e-008             wvth0=1.649609e-008              pvth0=-1.4115319e-014 k2=-0.0037834                 cit=0.00083648148              lcit=1.4688869e-009 voff=-0.12941025                lvoff=-2.4042266e-008            wvoff=-1.4274092e-008 pvoff=1.142648e-014              u0=0.055374619                lu0=6.3544045e-009 ua=-5.1003582e-011            lua=6.1300191e-017             wua=-4.1813745e-017 pua=2.0595971e-023             ub=3.8914728e-018             lub=-7.3851714e-025 wub=-1.7303361e-025            pub=1.5278868e-031             uc=-1.3968049e-011 luc=3.5644988e-017             wuc=1.8094305e-018             puc=-1.6254114e-023 vsat=191466.78                  lvsat=0.034613503                wvsat=-0.057730123 pvsat=2.6548387e-008             a0=19.208177                  la0=-1.0272154e-005 wa0=-2.0332248e-006            pa0=1.6145754e-012             ags=1.1477351 lags=2.9754388e-006             wags=1.2496066e-007             pags=-9.6653276e-014 keta=0.0088468588               lketa=-2.6717542e-008            wketa=-2.9064029e-008 pketa=-8.7484384e-015            pclm=1.1898096                  lpclm=9.8984042e-007 wpclm=5.5217788e-008             ppclm=-4.9602139e-013            pdiblc2=-0.020440362 lpdiblc2=7.102884e-008              wpdiblc2=2.4543774e-008             ppdiblc2=-2.1672153e-014 aigbacc=0.0094569283               laigbacc=1.5391323e-009             waigbacc=9.0811964e-010 paigbacc=-8.0186964e-016            aigc=0.011624397                laigc=-2.6698761e-010 waigc=-4.6247929e-011            paigc=3.9013667e-017             aigsd=0.0085207495 laigsd=3.548775e-010              waigsd=3.8517419e-012             paigsd=2.3384252e-019 tvoff=0.00725252                 ltvoff=-3.7483e-009               wtvoff=-1.86998e-009 ptvoff=1.65244e-015               kt1=-0.14655237                lkt1=-1.098139e-007 wkt1=-7.9248163e-008            pkt1=6.0015901e-014             kt2=-0.011505734 lkt2=-4.0806712e-009            wkt2=-1.96739e-009              pkt2=2.7627213e-015 ute=-2.0900586                 lute=1.7072963e-006             wute=2.523854e-008 pute=-2.2671781e-013            ua1=4.3654348e-009             lua1=-1.1556821e-015 wua1=-6.0699265e-016            pua1=1.3894066e-021             ub1=-1.3506428e-017 lub1=1.5289258e-023             wub1=3.5375011e-024             pub1=-5.6445121e-030 uc1=1.6224961e-010             luc1=-1.0445418e-018            wuc1=-9.3349948e-017 puc1=4.3344305e-023             at=78006.658                  pat=-8.1260726e-08 wat=0.009035997                lat=0.19778612                 wu0=0 pu0=0                          lk2=0                          wk2=0 pk2=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na_mac.8 nmos ( level=54                         lmin=4.5e-007                   lmax=9e-007 wmin=4.5e-07                    wmax=5.4e-007                   vth0=-0.059138324 lvth0=4.0202181e-008             wvth0=1.9424227e-008             pvth0=-1.6700865e-014 k2=-0.0015324088              lk2=-1.9876253e-009            wk2=-1.026452e-009 pk2=9.0635712e-016             cit=0.0023075556               lcit=1.6992844e-010 voff=-0.10810738                lvoff=-4.2852703e-008            wvoff=-1.8788046e-008 pvoff=1.5412302e-014             u0=0.05288311                 lu0=8.5544075e-009 wu0=3.544298e-009              pu0=-3.1296151e-015            ua=2.5803544e-010 lua=-2.1158126e-016            wua=-4.0741735e-017            pua=1.9649385e-023 ub=2.9679227e-018             lub=7.6977585e-026             wub=6.3885397e-026 pub=-5.6410806e-032            uc=8.285037e-011              luc=-4.9845677e-017 wuc=-4.3217316e-017            puc=2.3504502e-023             vsat=303795.56 lvsat=-0.064572809               wvsat=-0.067592373               pvsat=3.5256754e-008 a0=14.99427                   la0=-6.551274e-006             wa0=-2.7691799e-006 pa0=2.2644238e-012             ags=0.30755302                 lags=3.7173196e-006 wags=6.767228e-007              pags=-5.8385924e-013            keta=-0.060717321 lketa=3.4707629e-008             wketa=-2.2331314e-008            pketa=-1.4693426e-014 pclm=0.77474718                 lpclm=1.3563405e-006             wpclm=2.7074449e-007 ppclm=-6.8633147e-013            pdiblc2=0.097335505                lpdiblc2=-3.2967251e-008 wpdiblc2=-1.9218857e-008            ppdiblc2=1.6970251e-014             aigbacc=0.0112 aigc=0.011533197                laigc=-1.8645859e-010            waigc=-5.3553277e-011 paigc=4.5464289e-017             aigsd=0.0087758735               laigsd=1.2960293e-010 waigsd=4.0724883e-012             paigsd=3.8923456e-020             tvoff=0.00225952 ltvoff=6.60517e-010               wtvoff=4.88263e-010               ptvoff=-4.2989e-016 kt1=-0.34067339                lkt1=6.1594962e-008             wkt1=2.8049119e-008 pkt1=-3.4727599e-014            kt2=-0.012383073               lkt2=-3.3059813e-009 wkt2=-4.2245077e-011            pkt2=1.0628184e-015             ute=-0.15654067 wute=-2.3152002e-007            ua1=-1.2278344e-009            lua1=3.7831746e-015 wua1=3.6402532e-015             pua1=-2.3609114e-021            ub1=1.4615996e-017 lub1=-9.5428427e-024            wub1=-8.6685492e-024            pub1=5.1334303e-030 uc1=2.3252193e-010             luc1=-6.3094998e-017            wuc1=-8.6852665e-017 puc1=3.7607204e-023             at=569810.91                  lat=-0.23647704 wat=-0.17970711                pat=8.5399445e-08 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na_mac.9 nmos ( level=54                         lmin=2.7e-07                    lmax=4.5e-007 wmin=4.5e-07                    wmax=5.4e-007                   vth0=0.19265495 lvth0=-6.8824306e-008            wvth0=-1.0473667e-007            pvth0=3.7060804e-014 k2=-0.014895281               lk2=3.7984983e-009             wk2=5.0670176e-009 pk2=-1.7321152e-015            cit=-0.010512222               lcit=5.7208922e-009 wcit=5.8324933e-009             pcit=-2.5254696e-015            voff=-0.26713284 lvoff=2.6005323e-08              wvoff=7.0556386e-08              pvoff=-2.3273837e-14 u0=0.077296484                lu0=-2.0165837e-009            wu0=-2.5625752e-009 pu0=-4.85339e-016              ua=-1.0520847e-010            lua=-5.4296651e-017 wua=1.2106324e-016             pua=-5.0412168e-023            ub=2.7285124e-018 lub=1.8064224e-025             wub=4.7680595e-025             pub=-2.352054e-031 uc=-4.9508148e-011            luc=7.4655615e-018             wuc=2.6618916e-017 puc=-6.7345856e-024            vsat=160187.69                  lvsat=-0.0023906026 wvsat=0.0017004139               pvsat=5.2529768e-009             a0=-30.778472 la0=1.3268323e-005             wa0=1.9163919e-005             pa0=-7.2326082e-012 ags=25.795685                  lags=-7.3190417e-006            wags=-9.3924259e-006 pags=3.7760822e-012             keta=0.10754503                 lketa=-3.8149969e-008 wketa=-1.3417989e-007            pketa=3.3737007e-014             pclm=9.6987744 lpclm=-2.5077632e-006            wpclm=-3.9393275e-006            ppclm=1.1366297e-012 pdiblc2=0.0075160518               lpdiblc2=5.9245722e-009             wpdiblc2=4.4158814e-008 ppdiblc2=-1.0472281e-014            aigbacc=0.005757389                laigbacc=2.3566505e-009 waigbacc=3.7452384e-009             paigbacc=-1.6216882e-015            aigc=0.010991277 laigc=4.8193052e-011             waigc=1.8202994e-010             paigc=-5.6543244e-017 aigsd=0.0090749357               laigsd=1.0901586e-013             waigsd=4.3084264e-012 paigsd=-6.3237759e-020            tvoff=0.00396208                 ltvoff=-7.66908e-011 wtvoff=-1.96347e-010              ptvoff=-1.33454e-016              kt1=0.038827469 lkt1=-1.0272891e-007            wkt1=-1.5921897e-007            pkt1=4.6359485e-014 kt2=-0.03419288                lkt2=6.1376653e-009             wkt2=9.6912525e-009 pkt2=-3.1517861e-015            ute=-0.55805448                lute=1.7385548e-007 wute=2.1303263e-007             pute=-1.9249129e-013            ua1=6.0167507e-009 lua1=6.4626924e-016             wua1=-1.4425757e-015            pua1=-1.600465e-022 ub1=-8.7729299e-018            lub1=5.8456239e-025             wub1=6.5053258e-024 pub1=-1.4368575e-030            uc1=8.5352656e-011             luc1=6.2929814e-019 wuc1=4.8992944e-017             puc1=-2.1213945e-023            at=-210389.47 lat=0.10134973                 wat=0.19451009                 pat=-7.66366e-08 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_na12_mac.global nmos ( modelid=14                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 rdsmod=0                          igcmod=1                          igbmod=1 capmod=2                          rgatemod='1*rgflag_na12'            rbodymod=0 trnqsmod=0                          acnqsmod=0                          fnoimod=1.000000e+00 tnoimod=0.000000e+00               diomod=1                          tempmod=0 permod=1                          epsrox=3.9                        toxe=2.43e-009 toxm=2.43e-009                  dtox=2.15e-010                  xj=6.7e-008 ndep=1e+017                     ngate=3e+021                     nsd=1e+020 rsh=18.0                       rshg=16.42                      wint=0 lint=0                          dlc=1.2924e-008                dwc=0 xl=-1.2e-008                  xw=6e-009                     wl=0 wln=1                          ww=0                          wwn=1 wwl=0                          ll=0                          lln=1 lw=0                          lwn=1                          lwl=0 llc=0                          lwc=0                          lwlc=0 wlc=0                          wwc=0                          wwlc=0 phin=0.15                       k1=0.05                       k3=6.7881 k3b=0.456                      w0=0                          lpe0=5.5369e-006 lpeb=1e-008                     dvt0=0.000645                   dvt1=0.0021726 dvt2=0.1624                     dvtp0=1.1e-006                   dvtp1=3 dvt0w=0                          dvt1w=0                          dvt2w=0 ud=0                          b0=0                          b1=0 a1=0                          a2=1                          dwg=0 dwb=0                          voffl=0                          nfactor=1 eta0=0.02                       dsub=0.18                       cdsc=0 cdscb=0                          cdscd=0                          pclm=1.95 pdiblc1=0                          pdiblcb=1                          drout=0.56 pscbe1=1e+009                     pscbe2=1e-020                     pvag=1.5 delta=0.01                       fprout=300                        pdits=0.14 pditsl=0                          pditsd=0.37                       rdsw=120 prwg=0                          prwb=0                          wr=1 alpha0=0                          alpha1=0.0793                     beta0=10.75 bgidl=4.3391e+009                cgidl=0.295                      egidl=-0.3 cigbacc=0.11236                    nigbacc=3.7                        aigbinv=0.02 bigbinv=2e-005                     cigbinv=0.006                      eigbinv=1.1 nigbinv=1                          cigc=1.515e-005                 cigsd=0.015 dlcig=2.5e-009                   nigc=3.083                      poxedge=1 pigcd=3.3025                     ntox=1                          toxref=3e-009 vfbsdoff=0                          tnom=25                         kt1l=0 prt=0                          njs=1.02                       njd=1.02 xtis=3                          xtid=3                          tpb=0.0023 tpbsw=0.0018                     tpbswg=0.00252                    tcj=0.0023 tcjsw=0.00025                    tcjswg=0.00189                    tvfbsdoff=0.01015 xpart=1                          cgso=1.7433e-010                cgdo=1.7433e-010 cgbo=0                          cgsl=4e-011                     cgdl=4e-011 ckappas=0.6                        ckappad=0.6                        cf='6.7e-11+9.3e-11*ccoflag_na12' clc=0                          cle=0.6                        noff=3.7 voffcv=-0.29595                   acde=0.301                      moin=11.412 ijthsrev=0.01                       ijthdrev=0.01                       ijthsfwd=0.01 ijthdfwd=0.01                       xjbvs=1                          xjbvd=1 bvs=16.56                      bvd=16.56                      jss=1.28e-06 jsd=1.28e-06                   jsws=1.24e-12                   jswd=1.24e-12 jswgs=1.24e-12                   jswgd=1.24e-12                   jtsswgs=1e-010 jtsswgd=1e-010                     njtsswg=7                          xtsswgs=0.73768 xtsswgd=0.73768                    vtsswgs=2                          vtsswgd=2 tnjtsswg=1                          cjs=0.0001576                  cjd=0.0001576 mjs=0.34                       mjd=0.34                       mjsws=0.045 mjswd=0.045                      cjsws=2.102e-010                 cjswd=2.102e-010 cjswgs=1.551e-010                 cjswgd=1.551e-010                 mjswgs=0.479 mjswgd=0.479                      pbs=0.542                      pbd=0.542 pbsws=0.463                      pbswd=0.463                      pbswgs=0.881 pbswgd=0.881                      noia=0                          noib=0 noic=0                          em=1.000000e+06               ef=8.200000e-01 lintnoi=-1.300000e-07              dmcg=4.2e-008                   dmci=4.2e-008 dmdg=0                          dmcgt=0                          dwj=0 xgw=0                          xgl=2.64e-09                   ngcon=1 xrcrg1=12                         xrcrg2=1                          rbpb=50 rbpd=50                         rbps=50                         rbdb=50 rbsb=50                         gbmin=1e-012                     lpclm=0 ppclm=0                          weta0=0                          wpclm=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.11 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.62 sigma_factor='sigma_factor_na12' ccoflag='ccoflag_na12' rcoflag='rcoflag_na12' rgflag='rgflag_na12' mismatchflag='mismatchflag_mos_na12' globalflag='globalflag_mos_na12' totalflag='totalflag_mos_na12' global_factor='global_factor_na12' local_factor='local_factor_na12' sigma_factor_flicker='sigma_factor_flicker_na12' noiseflag='noiseflagn_na12' noiseflag_mc='noiseflagn_na12_mc' delvto=0 mulu0=1 dlc_fmt=2 par1='par1' par2='par2' par3='par3' par4='par4' par5='par5' par6='par6' par7='par7' par8='par8' par9='par9' par10='par10' par11='par11' par12='par12' par13='par13' par14='par14' par15='par15' par16='par16' par17='par17' par18='par18' par19='par19' par20='par20' par21='par21' par22='par22' par23='par23' par24='par24' par25='par25' par26='par26' par27='par27' par28='par28' par29='par29' par30='par30' par31='par31' par32='par32' w1='2.3875*0.35355' w2='0.70711*-0.35355' w3='0.54772*-0.0052117' w4='0.54772*-0.40307' w5='0.54772*-0.64548' w6='0.54772*-0.049915' w7='0.54772*-0.11513' w8='0.54772*-0.39385' w9='0' w10='0' tox_c='toxn_na12'                dxl_c='dxln_na12'                dxw_c='dxwn_na12' cgo_c='cgon_na12'                cgl_c='cgln_na12'                ddlc_c='ddlcn_na12' cj_c='cjn_na12'                 cjsw_c='cjswn_na12'               cjswg_c='cjswgn_na12' cf_c='cfn_na12'                 dvth_c='dvthn_na12'               dlvth_c='dlvthn_na12' dwvth_c='dwvthn_na12'              dpvth_c='dpvthn_na12'              du0_c='du0n_na12' dlu0_c='dlu0n_na12'               dwu0_c='dwu0n_na12'               dpu0_c='dpu0n_na12' dvsat_c='dvsatn_na12'              dwvsat_c='dwvsatn_na12'             dk2_c='dk2n_na12' dlk2_c='dlk2n_na12'               dwk2_c='dwk2n_na12'               dpk2_c='dpk2n_na12' deta0_c='deta0n_na12'              dweta0_c='dweta0n_na12'             dags_c='dagsn_na12' dlags_c='dlagsn_na12'              dwags_c='dwagsn_na12'              dpags_c='dpagsn_na12' dvoff_c='dvoffn_na12'              dlvoff_c='dlvoffn_na12'             dwvoff_c='dwvoffn_na12' dpvoff_c='dpvoffn_na12'             dcit_c='dcitn_na12'               dlcit_c='dlcitn_na12' dwcit_c='dwcitn_na12'              dpcit_c='dpcitn_na12'              dua_c='duan_na12' dlua_c='dluan_na12'               dwua_c='dwuan_na12'               dpua_c='dpuan_na12' dub_c='dubn_na12'                dlub_c='dlubn_na12'               dwub_c='dwubn_na12' dpub_c='dpubn_na12'               dkt1_c='dkt1n_na12'               dlkt1_c='dlkt1n_na12' dwkt1_c='dwkt1n_na12'              dpkt1_c='dpkt1n_na12'              dat_c='datn_na12' dlat_c='dlatn_na12'               dwat_c='dwatn_na12'               dpat_c='dpatn_na12' dpdiblc2_c='dpdiblc2n_na12'           dlpdiblc2_c='dlpdiblc2n_na12'          dwpdiblc2_c='dwpdiblc2n_na12' dppdiblc2_c='dppdiblc2n_na12'          dlvsat_c='dlvsatn_na12'             dpvsat_c='dpvsatn_na12' da0_c='da0n_na12'                dla0_c='dla0n_na12'               dwa0_c='dwa0n_na12' dpa0_c='dpa0n_na12'               ntox_c='ntoxn_na12'               dpclm_c='dpclmn_na12' dlpclm_c='dlpclmn_na12'             dwpclm_c='dwpclmn_na12'             dppclm_c='dppclmn_na12' duc1_c='duc1n_na12'               dluc1_c='dluc1n_na12'              dwuc1_c='dwuc1n_na12' dpuc1_c='dpuc1n_na12'              ff_flag_c='ff_flagn_na12'            monte_flag_c='monte_flagn_na12' c1f_c='c1fn_na12'                c2f_c='c2fn_na12'                c3f_c='c3fn_na12' global_mc='global_mc_flag_na12' tox_g='toxn_na12_ms_global'      dxl_g='dxln_na12_ms_global'      dxw_g='dxwn_na12_ms_global' cgo_g='cgon_na12_ms_global'      cgl_g='cgln_na12_ms_global'      cj_g='cjn_na12_ms_global' cjsw_g='cjswn_na12_ms_global'     cjswg_g='cjswgn_na12_ms_global' cf_g='cfn_na12_ms_global'       dvth_g='dvthn_na12_ms_global' dlvth_g='dlvthn_na12_ms_global'    dwvth_g='dwvthn_na12_ms_global' dpvth_g='dpvthn_na12_ms_global'    du0_g='du0n_na12_ms_global' dlu0_g='dlu0n_na12_ms_global'     dwu0_g='dwu0n_na12_ms_global' dpu0_g='dpu0n_na12_ms_global'     dvsat_g='dvsatn_na12_ms_global' dwvsat_g='dwvsatn_na12_ms_global'   dk2_g='dk2n_na12_ms_global' dlk2_g='dlk2n_na12_ms_global'     dweta0_g='dweta0n_na12_ms_global' dlcit_g='dlcitn_na12_ms_global'    dpcit_g='dpcitn_na12_ms_global' dat_g='datn_na12_ms_global'      dlat_g='dlatn_na12_ms_global' dwat_g='dwatn_na12_ms_global'     dpat_g='dpatn_na12_ms_global' dppdiblc2_g='dppdiblc2n_na12_ms_global'                                        dlvsat_g='dlvsatn_na12_ms_global' dpvsat_g='dpvsatn_na12_ms_global'   ntox_g='ntoxn_na12_ms_global' dpclm_g='dpclmn_na12_ms_global'    dwpclm_g='dwpclmn_na12_ms_global' dppclm_g='dppclmn_na12_ms_global'   ff_flag_g='ff_flagn_na12_ms_global' monte_flag_g='monte_flagn_na12_ms_global'                                      ddlc_g='ddlcn_na12_ms_global' dpdiblc2_g='dpdiblc2n_na12_ms_global' weight1=-3.3429333 weight2=1.6658 weight3=1.5021333 weight4=0.66666667 weight5=-0.45894667 tox_1=4.5171226e-012 tox_2=1.7501088e-012 tox_3=-1.3078065e-011 tox_4=-3.7477187e-011 tox_5=2.2526113e-012 dxl_1=2.2159111e-010 dxl_2=8.5853429e-011 dxl_3=-6.4155321e-010 dxl_4=1.8385092e-009 dxl_5=1.1050055e-010 dxw_1=-6.8569343e-010 dxw_2=2.6888134e-011 dxw_3=-1.2625063e-009 dxw_4=-1.3829069e-024 dxw_5=-5.8250291e-009 cgo_1=-1.2035e-012 cgo_2=-1.7632e-013 cgo_3=3.481e-013 cgo_4=-6.8407e-028 cgo_5=6.6695e-014 cgl_1=-2.7613e-013 cgl_2=-4.0457e-014 cgl_3=7.9872e-014 cgl_4=-8.5995e-029 cgl_5=1.5303e-014 cj_1=1.088e-006 cj_2=1.594e-007 cj_3=-3.147e-007 cj_4=2.6238e-021 cj_5=-6.0295e-008 cjsw_1=1.4511e-012 cjsw_2=2.126e-013 cjsw_3=-4.1973e-013 cjsw_4=1.0126e-027 cjsw_5=-8.0418e-014 cjswg_1=1.0707e-012 cjswg_2=1.5687e-013 cjswg_3=-3.097e-013 cjswg_4=1.332e-028 cjswg_5=-5.9338e-014 cf_1=-4.6252e-013 cf_2=-6.7765e-014 cf_3=1.3379e-013 cf_4=-5.6362e-028 cf_5=2.5633e-014 dvth_1=0.0043417 dvth_2=0.00032499 dvth_3=0.0020537 dvth_4=-9.2266e-019 dvth_5=-0.00094626 dlvth_1=1.4054e-009 dlvth_2=1.5804e-011 dlvth_3=7.7215e-010 dlvth_4=-1.0534e-024 dlvth_5=-3.259e-010 dwvth_1=1.6591e-009 dwvth_2=-4.4071e-011 dwvth_3=7.6516e-010 dwvth_4=-7.3399e-024 dwvth_5=-3.5519e-010 dpvth_1=1.5717e-016 dpvth_2=-2.8981e-016 dpvth_3=1.8065e-016 dpvth_4=-9.4455e-031 dpvth_5=-5.7372e-017 du0_1=0.00027684 du0_2=-5.445e-005 du0_3=0.00065658 du0_4=2.0208e-019 du0_5=-0.00018549 dlu0_1=7.4972e-011 dlu0_2=-1.0615e-011 dlu0_3=1.5624e-010 dlu0_4=5.8462e-026 dlu0_5=-4.3936e-011 dwu0_1=9.494e-011 dwu0_2=-5.0265e-013 dwu0_3=7.2728e-011 dwu0_4=6.3728e-026 dwu0_5=-2.8514e-011 dpu0_1=-3.0256e-017 dpu0_2=-3.6254e-017 dpu0_3=9.0108e-017 dpu0_4=1.4976e-031 dpu0_5=-1.7158e-017 dvsat_1=754.47 dvsat_2=88.179 dvsat_3=882.03 dvsat_4=1.7536e-012 dvsat_5=-245.73 dwvsat_1=0.0002455 dwvsat_2=0.00026283 dwvsat_3=0.0010909 dwvsat_4=2.2808e-019 dwvsat_5=-0.00026071 dk2_1=3.1151e-005 dk2_2=-4.8239e-005 dk2_3=-1.4528e-005 dk2_4=7.7589e-020 dk2_5=-7.4777e-007 dlk2_1=7.7851e-011 dlk2_2=4.6608e-011 dlk2_3=-1.8841e-011 dlk2_4=9.2358e-026 dlk2_5=-4.9669e-012 dweta0_1=1.868e-010 dweta0_2=3.7939e-010 dweta0_3=-1.725e-011 dweta0_4=1.0046e-025 dweta0_5=-1.6877e-011 dlcit_1=-5.1918e-012 dlcit_2=8.0399e-012 dlcit_3=2.4213e-012 dlcit_4=-2.0267e-026 dlcit_5=1.2463e-013 dpcit_1=4.67e-018 dpcit_2=9.4848e-018 dpcit_3=-4.3126e-019 dpcit_4=-1.0724e-032 dpcit_5=-4.2191e-019 dat_1=2995 dat_2=42.774 dat_3=-907.68 dat_4=-1.6444e-011 dat_5=-158.64 dlat_1=-0.00036958 dlat_2=0.00010426 dlat_3=0.00012346 dlat_4=-1.7629e-019 dlat_5=1.7547e-005 dwat_1=0.00020767 dwat_2=-0.0003216 dwat_3=-9.6853e-005 dwat_4=3.1086e-019 dwat_5=-4.9852e-006 dpat_1=-1.0384e-010 dpat_2=1.608e-010 dpat_3=4.8426e-011 dpat_4=-4.3198e-025 dpat_5=2.4926e-012 dppdiblc2_1=-5.1918e-017 dppdiblc2_2=8.0399e-017 dppdiblc2_3=2.4213e-017 dppdiblc2_4=3.4659e-032 dppdiblc2_5=1.2463e-018 dlvsat_1=0.00017644 dlvsat_2=0.00022826 dlvsat_3=-2.9887e-005 dlvsat_4=-1.3123e-019 dlvsat_5=-1.353e-005 dpvsat_1=1.0782e-010 dpvsat_2=-7.8369e-011 dpvsat_3=-4.1027e-011 dpvsat_4=-2.0889e-025 dpvsat_5=-4.2302e-012 ntox_1=-0.13702 ntox_2=-0.055278 ntox_3=0.035956 ntox_4=4.2145e-016 ntox_5=0.0082462 dpclm_1=-0.01868 dpclm_2=-0.037939 dpclm_3=0.001725 dpclm_4=-4.1205e-018 dpclm_5=0.0016877 dwpclm_1=-4.67e-009 dwpclm_2=-9.4848e-009 dwpclm_3=4.3126e-010 dwpclm_4=-1.3466e-023 dwpclm_5=4.2191e-010 dppclm_1=2.1669e-015 dppclm_2=4.4009e-015 dppclm_3=-2.0011e-016 dppclm_4=5.3959e-030 dppclm_5=-1.9577e-016 ff_flag_1=-0.051918 ff_flag_2=0.080399 ff_flag_3=0.024213 ff_flag_4=6.8785e-017 ff_flag_5=0.0012463 monte_flag_1=0.0852269 monte_flag_2=0.0330204 monte_flag_3=-0.24675 monte_flag_4=0.707115 monte_flag_5=0.0425 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.992854610120824 b_4=0.00136015580096095        c_4=-0.0170970888345293        d_4=0.00322840519628978 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=0                          g_4_2=0 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1='0.0085-0.0007'            mis_a_2=0.55                       mis_a_3=0 mis_b_1='0.003-0.001'              mis_b_2=0                          mis_b_3=0 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.0038                     mis_d_2=0                          mis_d_3=0 mis_e_1=0.026                      mis_e_2='0.5+0.01'                 mis_e_3=0 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=6e-09                      xl0=-1.2e-08 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18                         bidirectionflag=1 designflag=1 cf0=6.7e-11                    cco=9.3e-11 noimod=1                          noic2='2.236'                    noic3='0.6' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.453e-6            sbref0=0.453e-6 samax=10e-6		sbmax=10e-6 samin=0.072e-6            sbmin=0.072e-6 rllodflag=0                  lreflod=0.9e-6              llodref=1 lod_clamp=-1e90 wlod0=0 ku00=0                   lku00=0                   wku00=0 pku00=0                   tku00=0                   llodku00=1 wlodku00=1                   kvsat0=0 kvth00=-0e-9               lkvth00=0e-8                wkvth00=0e-8 pkvth00=0                   llodvth0=1                   wlodvth0=1 stk20=0                   lodk20=1                   steta00=0e-11 lodeta00=1 wlod00=0 ku000=-0e-9               lku000=0e-28               wku000=0         		pku000=0 llodku000=1                   wlodku000=1 kvth000=0.0e-8              lkvth000=0e-23               wkvth000=-0e-16         	pkvth000=0 llodvth00=1                   wlodvth00=1                   steta000=0 stk200=0                   lodk200=1 lodeta000=1 wlod1=0                   llod1=1e-6 ku01=-2e-7               lku01=2.9e-19            wku01=0 pku01=0                   llodku01=2 wlodku01=1                   kvsat1=-2 kvth01=1.5e-7              lkvth01=-1.15e-13             wkvth01=0 pkvth01=0                   llodvth1=1                  wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=-0.00               lku02=0.0e-7              wku02=0 pku02=0                   tku02=0                   llodku02=1 wlodku02=1                   kvsat2=0 kvth02=0e-3               lkvth02=0e-7                   wkvth02=0 pkvth02=0                   llodvth2=1                   wlodvth2=1 stk22=0                   lodk22=1                   steta02=0e-4 lodeta02=1 wlod02=0 ku002=0             lku002=-0e-18              wku002=0e-9         		pku002=0 llodku002=1                   wlodku002=1 kvth002=0e-3                lkvth002=-0e-15               wkvth002=0e-9         	    pkvth002=0 llodvth02=2                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0.0                 lku03=0                   wku03=0 pku03=0                   tku03=0                   llodku03=1 wlodku03=1                   kvsat3=0.0 kvth03=0e-3                lkvth03=0                   wkvth03=0 pkvth03=0                   llodvth3=1                   wlodvth3=1 stk23=0                   lodk23=1                   steta03=0 lodeta03=1 wlod03=0 ku003=0                   lku003=0                   wku003=0e-9         		pku003=-0e-16 llodku003=1                   wlodku003=1 kvth003=0e-3                lkvth003=-0e-9               wkvth003=0e-10         	pkvth003=-0e-18 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=1.93e-7             sa_b1=0.99e-7             dpdbinflag=1 w_b=9e-6                w_b1=10e-6 sparef=1.54e-7             spamax=4.8e-7              spamin=1.54e-7 kvth0dpc=0                   wkvth0dpc=0e-7              wdpckvth0=1 lkvth0dpc=0e-8                ldpckvth0=1                 pkvth0dpc=0e-15 ku0dpc=0                   wku0dpc=0e-7              wdpcku0=1 lku0dpc=0e-7                ldpcku0=1                 pku0dpc=0e-14 keta0dpc=0                   wketa0dpc=0e-9              wdpcketa0=1 kvsatdpc=0                  wdpc=0 kvth0dpc_b1=0.00              kvth0dpc_b2=-0.000          dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=0.8                  wkvth0dpl=0e-7              wdplkvth0=1 lkvth0dpl=-0e-7               ldplkvth0=1                 pkvth0dpl=0.00e+00 ku0dpl=-0.5                   wku0dpl=0e-7                wdplku0=1 lku0dpl=0e-7                  ldplku0=1                   pku0dpl=0e-13 keta0dpl=0                    wketa0dpl=0.00e+00          wdplketa0=1 kvsatdpl=0                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000          dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=-0.0                wkvth0dpx=0e-6              wdpxkvth0=1 lkvth0dpx=0e-7                ldpxkvth0=1.0               pkvth0dpx=0e-14 ku0dpx=0.0                 wku0dpx=0e-6              wdpxku0=1 lku0dpx=0e-8                ldpxku0=1.0               pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7              wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000          dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=-0.025                  wkvth0dps=0                 wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0               pkvth0dps=0 ku0dps=-0                  wku0dps=-0.0e-9           wdpsku0=1 lku0dps=0.0e-16             ldpsku0=1.0               pku0dps=0.0e-23 keta0dps=0.00                wketa0dps=0                 wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000          dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=0.00                 wkvth0dpa=-0e-08            wdpakvth0=1 lkvth0dpa=0.00e+00            ldpakvth0=1                 pkvth0dpa=0.00e+00 ku0dpa=0.08                   wku0dpa=4e-9              wdpaku0=1 lku0dpa=-1e-08                ldpaku0=1                   pku0dpa=0.00e+00 keta0dpa=0                    wketa0dpa=0.00e+00          wdpaketa0=1 ka0dpa=0                      wka0dpa=0                   wdpaka0=1 lka0dpa=0.00e+00              ldpaka0=1                   pka0dpa=0.00e+00 kvsatdpa=0                    wdpa=0 kvth0dpa_b1=0.000             kvth0dpa_b2=-0.00           dpabinflg=0 ku0dpa_b1=-0.00             ku0dpa_b2=0.00 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.08e-7             spbmax='4.8e-7+6.8e-7'     spbmin='1.54e-7+3.54e-7' pse_mode=1 kvth0dp2=0              	 wkvth0dp2=0            		 wdp2kvth0=1 lkvth0dp2=0e-8           	 ldp2kvth0=1                   pkvth0dp2=0 ku0dp2=0            	     wku0dp2=0e-9             	 wdp2ku0=1 lku0dp2=0.0e-8          	 ldp2ku0=1                 	 pku0dp2=0 keta0dp2=0               	 wketa0dp2=0               	 wdp2keta0=1 kvsatdp2=0.0               	 wdp2=0 kvth0dp2l=1                  wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0e-8               ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0               wku0dp2l=0e-8               wdp2lku0=1 lku0dp2l=0e-8               ldp2lku0=1                  pku0dp2l=0e-15 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0.0                wdp2l=0 kvth0dp2l_b1=0.00             kvth0dp2l_b2=-0.00            dp2lbinflg=1 ku0dp2l_b1=0.0              ku0dp2l_b2=0.00 keta0dp2l_b1=0                keta0dp2l_b2=0 kvth0dp2a=0.0                wkvth0dp2a=0            		 wdp2akvth0=1 lkvth0dp2a=0e-9             	 ldp2akvth0=1                  pkvth0dp2a=0 ku0dp2a=-0.15               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=-0e-8              ldp2aku0=1                  pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1                  pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=0.0              kvth0dp2a_b2=0.0              dp2abinflg=0 ku0dp2a_b1=-0.0             ku0dp2a_b2=-0.0 keta0dp2a_b1=0                keta0dp2a_b2=0 ka0dp2a_b1=-0               ka0dp2a_b2=-0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1e-7 kvth0enx=-0.00            	 wkvth0enx=-0e-5             wenxkvth0=0.0 lkvth0enx=0          		 lenxkvth0=1                   pkvth0enx=-0.0e-12 ku0enx=-0         		 wku0enx=-0e-4      		 wenxku0=1 lku0enx=0e-8          	 lenxku0=1                   pku0enx=-0e-12 keta0enx=0.00                wketa0enx=0                   wenxketa0=1 ka0enx=0                   wka0enx=0                   wenxka0=1 lka0enx=0          		 lenxka0=1                   pka0enx=0 kvsatenx=0.0                 wenx=0                   ku0enx0=0 eny0=2e-6 enyref=2e-6             enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0.000          	 wkvth0eny=0       		     wenykvth0=1 lkvth0eny=0        			 lenykvth0=1                   pkvth0eny=0e-17 ku0eny=0          		 wku0eny=0e-8        		 wenyku0=1 ku0eny0=0.00          		 wku0eny0=0                   weny0ku0=1 lku0eny=0e-6       		 lenyku0=1                 	 pku0eny=0e-16 keta0eny=0               	 wketa0eny=0                   wenyketa0=1 ka0eny=0              	 wka0eny=0             		 wenyka0=1 lka0eny=0      		     lenyka0=1                	 pka0eny=0 kvsateny=0.0               	 weny=0 kvth0eny1=-0e-4          	 wkvth0eny1=0        		     weny1kvth0=1 lkvth0eny1=0             	 leny1kvth0=1                  pkvth0eny1=-0e-18 ku0eny1=-0.000        	 wku0eny1=-0e-9            	 weny1ku0=1 lku0eny1=0e-4      		 leny1ku0=0.0                pku0eny1=-0.0e-12 keta0eny1=0              	 wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1                	 pka0eny1=0 kvsateny1=0.0                weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.8126e-5           ringxmin=0 kvth0rx=0.00              	 wkvth0rx=0e-9          	     wrxkvth0=1 lkvth0rx=0              	 lrxkvth0=1                	 pkvth0rx=0e-16 ku0rx=0              	 wku0rx=0e-8           	 wrxku0=1 lku0rx=0e-9        		 lrxku0=1                   pku0rx=0 keta0rx=0                	 wketa0rx=0                   wrxketa0=1 kvsatrx=0.1                 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=1.6027e-5           ringymin=0 kvth0ry=-0.000           	 wkvth0ry=0           	     wrykvth0=1 lkvth0ry=0              	 lrykvth0=1                 	 pkvth0ry=0 ku0ry=-0.0          	 wku0ry=0           		 wryku0=1 lku0ry=0        			 lryku0=1                 	 pku0ry=0 keta0ry=0                	 wketa0ry=0                   wryketa0=1 kvsatry=0.0                 wry=0 kvth0ry0=0                	 ku0ry0=0 sfxref=8.26e-7           sfxmax=10e-6             minwodx=0.0e-6 sfxmin=0.252e-6 lrefodx=5e-8              lodxref=1                 wodx=0e-6 kvth0odxa=-0.000            lkvth0odxa=0.0e-13           lodxakvth0=2.0 wkvth0odxa=0.0e-7            wodxakvth0=1.0               pkvth0odxa=0.0e-16 ku0odxa=-0.00             lku0odxa=0.0e-13           lodxaku0=2.0 wku0odxa=0.0e-7            wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.00              wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a='-0.000'            lkvth0odx1a='1.0e-13*0'           lodx1akvth0='2.0' wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.90 kvth0odx1b=-0.0009           lkvth0odx1b='0+3e-12-1e-12'            lodx1bkvth0=1.0 wkvth0odx1b=-0.0e-5           wodx1bkvth0=1.0               pkvth0odx1b=0.0e-16 ku0odx1b='-0.0028-0.0005*3'           lku0odx1b='1.1e-10+0.5e-10'           lodx1bku0=1.0 wku0odx1b=-0.8e-10          wodx1bku0=1.0               pku0odx1b=0.0e-16 sfyref=7.92e-7 sfymin=0.15e-6 sfymax=10e-6             minwody=0.9e-6            wody=5e-7 kvth0odya=-0.00             lkvth0odya=0.0e-13           lodyakvth0=1.0 wkvth0odya=-0.0e-6           wodyakvth0=0.5               pkvth0odya=0.0e-16 ku0odya=-0.00             lku0odya=0.0e-13           lodyaku0=1.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=1.2 lrefody=5e-8              lodyref=1 kvth0odyb=0.018             lkvth0odyb=-8.0e-10          lodybkvth0=1.0 wkvth0odyb=-12.5e-8          wodybkvth0=1.0               pkvth0odyb=-0.5e-15 ku0odyb=0.01              lku0odyb=0.15e-8           lodybku0=1.0 wku0odyb=-0.5e-7           wodybku0=1.0               pku0odyb=0.2e-15 web_mac=0  wec_mac=0 kvsatwe=0 lodflag=1    pseflag=1 ceslflag=0 oseflag=1 wpeflag=0 )
.model nch_na12_mac.1 nmos ( lmin=9e-007                     lmax=9.019e-06                  wmin=9e-007 wmax=9.001e-06                  level=54                         vth0=0.04037136 lvth0=8.9294766e-009             wvth0=-2.6452478e-008            pvth0=2.3665126e-014 k2=-0.010425207               lk2=-3.6653923e-010            wk2=5.8102003e-009 pk2=-1.7127985e-015            u0=0.071819578                lu0=1.0292613e-009 wu0=-6.0347517e-009            pu0=1.1007728e-014             ua=1.3561181e-009 lua=-8.7930897e-016            wua=1.5955162e-016             pua=-4.8795302e-023 ub=2.0954958e-018             lub=6.2350668e-025             wub=-5.903862e-025 pub=6.8706484e-031             uc=-4.3437123e-011            luc=1.9524330e-017 wuc=5.4508554e-018             puc=-1.1364064e-023            vsat=127200 a0=4.8020385                  la0=4.3759236e-006             wa0=4.6928932e-006 pa0=-8.6520343e-012            ags=2.7898648                  lags=-1.8769588e-007 wags=-1.4090245e-006            pags=2.021392e-012              keta=-0.050476836 lketa=1.9352602e-008             wketa=-1.4636572e-008            pketa=-4.1380719e-015 voff=-0.09533977                lvoff=-2.5826875e-008            wvoff=-4.1804219e-010 pvoff=-1.0792338e-014            minv=-0.50904892                lminv=4.1850333e-007 wminv=6.6551285e-008             pminv=-3.9689360e-013            etab=-0.032316098 wetab=1.4185331e-008             cit=0.0026067601               lcit=4.0923792e-010 wcit=1.2775341e-010             pcit=4.4705866e-016             pdiblc2=0.020556292 lpdiblc2=2.5865226e-009             wpdiblc2=3.48846e-009               ppdiblc2=4.4993715e-015 agidl=2.3004085e-006             lagidl=1.6257308e-013             wagidl=6.1340021e-012 pagidl=-2.8005684e-018            aigbacc=0.013452136                laigbacc=4.8650361e-010 waigbacc=-6.2595223e-011            paigbacc=5.5584558e-017             bigbacc=0.0050672974 lbigbacc=-5.7972220e-011            wbigbacc=-6.0608007e-010            pbigbacc=5.2209782e-016 aigc=0.012412419                laigc=-1.6483337e-010            waigc=-2.0820211e-011 paigc=-1.7181187e-016            bigc=0.0015455                  aigsd=0.010040862 laigsd=2.6505353e-010             waigsd=-1.3003710e-010            paigsd=1.3669623e-016 bigsd=0.00043914521              lbigsd=2.0538451e-010             wbigsd=-1.0643779e-010 pbigsd=1.0703998e-016             ute=-1.6692422                 lute=4.7586736e-007 wute=4.6235073e-007             pute=-3.8373197e-013            kt1=-0.17468752 lkt1=-1.1676165e-007            wkt1=-1.8892598e-008            pkt1=5.4730938e-014 kt2=-0.013851892               lkt2=5.1042630e-009             wkt2=-1.0780792e-009 pkt2=-1.2383446e-015            ua1=3.9080069e-009             lua1=6.2097506e-016 wua1=9.8244266e-016             pua1=-5.0055880e-022            ub1=-6.2983503e-018 lub1=2.5127729e-024             wub1=1.5628923e-024             pub1=-2.1983693e-030 uc1=-4.2855099e-012            luc1=2.4669819e-017             wuc1=1.8848814e-017 puc1=-4.4694948e-023            at=101481.88                  lat=0.031431744 wat=6.5753041e-005             pat=-1.5077311e-008            tvoff=0.007075295 ltvoff=-5.3165864e-009            wtvoff=-1.2624097e-009            ptvoff=2.0155358e-015 lvsat=0                          wvsat=0                          pvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na12_mac.2 nmos ( lmin=4.5e-007                   lmax=9e-007                     wmin=9e-007 wmax=9.001e-06                  level=54                         vth0=0.045515233 lvth0=4.3617173e-009             wvth0=1.148271e-008              pvth0=-1.0021322e-014 k2=-0.0098942763              lk2=-8.3800568e-010            wk2=3.4557488e-009 pk2=3.7795446e-016             u0=0.066135746                lu0=6.0765038e-009 wu0=2.1433206e-008             pu0=-1.3383819e-014            ua=4.9222281e-010 lua=-1.1216994e-016            wua=4.7532462e-016             pua=-3.2920173e-022 ub=2.612555e-018              lub=1.6435807e-025             wub=8.0534909e-025 pub=-5.5234809e-031            uc=-3.0092693e-011            luc=7.6744765e-018 wuc=-8.9839084e-018            puc=1.4540059e-024             vsat=127200 a0=12.982329                  la0=-2.8881744e-006            wa0=-3.9490206e-006 pa0=-9.7801484e-013            ags=2.7089327                  lags=-1.1582816e-007 wags=1.7061146e-006             pags=-7.448515e-013             keta=-0.056262247 lketa=2.4490046e-008             wketa=-3.6430390e-008            pketa=1.5214839e-014 voff=-0.096425817               lvoff=-2.4862466e-008            wvoff=-3.435774e-008 pvoff=1.9346114e-014             minv=-0.036497415               lminv=-1.1224060e-009 wminv=-3.9178428e-007            pminv=1.0108388e-014             etab=-0.032316098 wetab=1.4185331e-008             cit=0.0047975495               lcit=-1.5361831e-009 wcit=-1.4693727e-009            pcit=1.8653067e-015             pdiblc2=0.031386592 lpdiblc2=-7.0307842e-009            wpdiblc2=8.3758927e-009             ppdiblc2=1.5933118e-016 agidl=1.2662283e-006             lagidl=1.0809251e-012             wagidl=4.2697301e-012 pagidl=-1.1450949e-018            aigbacc=0.014                      bigbacc=0.005003973 lbigbacc=-1.7401643e-012            wbigbacc=-3.5780638e-011            pbigbacc=1.5671919e-017 aigc=0.012367461                laigc=-1.2491133e-010            waigc=-2.9547169e-010 paigc=7.2078640e-017             bigc=0.0015455                  aigsd=0.010298432 laigsd=3.6331642e-011             waigsd=4.9267937e-011             paigsd=-2.2526643e-017 bigsd=0.00064165657              lbigsd=2.5554421e-011             wbigsd=2.7829385e-011 pbigsd=-1.2189271e-017            ute=-0.89319075                lute=-2.1326635e-007 wute=-2.8902536e-008            pute=5.2500930e-014             kt1=-0.33432739 lkt1=2.4998548e-008             wkt1=1.317391e-007              pkt1=-7.9030007e-014 kt2=-0.0043143254              lkt2=-3.3650965e-009            wkt2=-1.9006019e-009 pkt2=-5.0794432e-016            ua1=5.43933e-009               lua1=-7.3883982e-016 wua1=-8.1096064e-017            pua1=4.4386358e-022             ub1=-2.964041e-018 lub1=-4.4809371e-025            wub1=-7.2371310e-025            pub1=-1.6786367e-031 uc1=4.3388816e-011             luc1=-1.7664982e-017            wuc1=-3.5322877e-017 puc1=3.4095131e-024             at=247468.69                  lat=-0.098204542 wat=-0.060922822               pat=3.9080543e-008             tvoff=0.0010680198 ltvoff=1.7873946e-011             wtvoff=2.3483340e-009             ptvoff=-1.1908047e-015 lvsat=0                          wvsat=0                          pvsat=0 vsat_mc=380.995                    lvsat_mc=-0.000338324               wvsat_mc=-0.00343162 pvsat_mc=3.04728e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na12_mac.3 nmos ( lmin=2.7e-07                    lmax=4.5e-007                   wmin=9e-007 wmax=9.001e-06                  level=54                         vth0=0.038145261 lvth0=7.5897653e-009             wvth0=1.051486e-008              pvth0=-9.5974034e-015 k2=-0.016792483               lk2=2.183409e-009              wk2=5.4581456e-009 pk2=-4.9909533e-016            u0=0.093295559                lu0=-5.8194944e-009 wu0=-1.4747257e-008            pu0=2.4632239e-015             ua=1.3312289e-009 lua=-4.7965462e-016            wua=-6.1544527e-016            pua=1.4855549e-022 ub=2.9532418e-018             lub=1.5137281e-026             wub=-5.8465549e-025 pub=5.6473914e-032             uc=-3.0466867e-011            luc=7.8383648e-018 wuc=-2.6880204e-017            puc=9.2925834e-024             vsat=152513.96 a0=13.758751                  la0=-3.2282473e-006            wa0=-1.732023e-005 pa0=4.8785747e-012             ags=3.7671741                  lags=-5.7933789e-007 wags=3.1784529e-007             pags=-1.3678956e-013            keta=-0.024168945 lketa=1.0433180e-008             wketa=-8.9645185e-009            pketa=3.1847873e-015 voff=-0.14573641                lvoff=-3.2644251e-009            wvoff=1.2395963e-008 pvoff=-1.1320079e-015            minv=-0.086153322               lminv=2.0626881e-008 wminv=-8.0135278e-007            pminv=1.8949939e-013             etab=-0.055869106 wetab=2.0050108e-008             cit=-0.0019865447              lcit=1.4352502e-009 wcit=8.2091011e-009             pcit=-2.3738649e-015            pdiblc2=0.015452665 lpdiblc2=-5.1724209e-011            wpdiblc2=2.3140631e-008             ppdiblc2=-6.307624e-015 agidl=1.6960081e-006             lagidl=8.9268156e-013             wagidl=2.1280749e-012 pagidl=-2.0704994e-019            aigbacc=0.014022445                laigbacc=-9.8308830e-012 waigbacc=-2.0213911e-010            paigbacc=8.8536932e-017             bigbacc=0.005 aigc=0.012254957                laigc=-7.5634402e-011            waigc=-1.8414769e-010 paigc=2.3318731e-017             bigc=0.0015455                  aigsd=0.010385448 laigsd=-1.7811542e-012            waigsd=-1.2607571e-011            paigsd=4.5748298e-018 bigsd=0.0007                     ute=-1.953402                  lute=2.5110617e-007 wute=1.6929151e-007             pute=-3.4308061e-014            kt1=-0.3023336 lkt1=1.0985268e-008             wkt1=-1.1532842e-007            pkt1=2.9185567e-014 kt2=-0.018407434               lkt2=2.8076853e-009             wkt2=2.4292286e-009 pkt2=-2.4044101e-015            ua1=3.6347668e-009             lua1=5.1558889e-017 wua1=2.5862222e-015             pua1=-7.2442183e-022            ub1=-5.8376224e-018 lub1=8.1053496e-025             wub1=-2.8293331e-024            pub1=7.5439790e-031 uc1=-1.8788085e-012            luc1=2.1622371e-018             wuc1=-5.020417e-017 puc1=9.9275197e-024             at=-3997.0928                 lat=0.011937472 wat=0.059473457                pat=-1.3653027e-008            tvoff=0.00071577756 ltvoff=1.7215606e-010             wtvoff=-1.1304412e-009            ptvoff=3.3289886e-016 lvsat=-0.011087515               wvsat=0.0025700545               pvsat=-1.1256838e-009 letab=1.0316217e-008             petab=-2.5687726e-015            vth0_mc=0.00573334 lvth0_mc=-2.5112e-09                wvth0_mc=1.5e-15                    pvth0_mc=4.8e-21 vsat_mc=3427.66                    lvsat_mc=-0.00167277                wvsat_mc=0.00785714 pvsat_mc=-1.89719e-09 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na12_mac.4 nmos ( lmin=9e-007                     lmax=9.019e-06                  wmin=5.4e-007 wmax=9e-007                     level=54                         vth0=0.0049139464 lvth0=6.7135748e-008             wvth0=5.6719387e-009             pvth0=-2.9069757e-014 k2=-0.012588084               lk2=1.8044193e-009             wk2=7.7697666e-009 pk2=-3.6796869e-015            u0=0.070237351                lu0=3.1451701e-008 wu0=-4.6012543e-009            pu0=-1.6555003e-014            ua=1.7238973e-009 lua=-5.6617503e-016            wua=-1.7365636e-016            pua=-3.3249465e-022 ub=2.2955323e-018             lub=1.5843543e-024             wub=-7.7161924e-025 pub=-1.8346307e-031            uc=-2.7643688e-011            luc=-1.1351409e-018 wuc=-8.8579962e-018            puc=7.3534163e-024             vsat=127200 a0=10.093339                  la0=-4.9286934e-006            wa0=-1.0102485e-007 pa0=-2.2205124e-013            ags=1.4085497                  lags=2.842802e-006 wags=-1.5755308e-007            pags=-7.2423907e-013            keta=-0.079695973 lketa=2.8289036e-008             wketa=1.1835966e-008             pketa=-1.2234482e-014 voff=-0.095126662               lvoff=-7.1065164e-008            wvoff=-6.1111825e-010 pvoff=3.0193552e-014             minv=-0.40314887                lminv=-4.7126716e-008 wminv=-2.9394157e-008            pminv=2.4967225e-014             etab=-0.033219332 wetab=1.5003660e-008             cit=0.00074651113              lcit=2.338248e-009 wcit=1.813139e-009              pcit=-1.3006245e-015            pdiblc2=0.030188198 lpdiblc2=1.1683374e-008             wpdiblc2=-5.2380468e-009            ppdiblc2=-3.7423757e-015 agidl=1.691855e-005              lagidl=-5.0139856e-011            wagidl=-7.1100339e-012 pagidl=4.2773432e-017             aigbacc=0.013807793                laigbacc=6.0165539e-010 waigbacc=-3.8482129e-010            paigbacc=-4.8742955e-017            bigbacc=0.0050204647 lbigbacc=3.7931091e-010             wbigbacc=-5.6364971e-010            pbigbacc=1.2591930e-016 aigc=0.012639971                laigc=-5.6312768e-010            waigc=-2.2698291e-010 paigc=1.8904278e-016             bigc=0.0015455                  aigsd=0.010034415 laigsd=2.6975432e-010             waigsd=-1.2419571e-010            paigsd=1.3243732e-016 bigsd=0.00042991614              lbigsd=2.0854726e-010             wbigsd=-9.8076255e-011 pbigsd=1.0417453e-016             ute=-0.71514534                lute=-2.8437726e-007 wute=-4.0206105e-007            pute=3.0504966e-013             kt1=-0.25867339 lkt1=-8.828746e-009             wkt1=5.7198592e-008             pkt1=-4.3056277e-014 kt2=-0.003752336               lkt2=-3.9320765e-009            wkt2=-1.0228277e-008 pkt2=6.9485790e-015             ua1=8.2610491e-009             lua1=-1.5014370e-015 wua1=-2.9614135e-015            pua1=1.4223465e-021             ub1=-5.9634497e-018 lub1=1.0593526e-024             wub1=1.2594724e-024             pub1=-8.8157049e-031 uc1=1.9153891e-011             luc1=-3.0197399e-018            wuc1=-2.387284e-018 puc1=-1.9608207e-023            at=101986.72                  lat=0.0119955 wat=-0.00039162868             pat=2.5319257e-009             tvoff=0.0019057486 ltvoff=-1.3514977e-009            wtvoff=3.4211994e-009             ptvoff=-1.5768346e-015 lvsat=0                          wvsat=0                          pvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na12_mac.5 nmos ( lmin=4.5e-007                   lmax=9e-007                     wmin=5.4e-007 wmax=9e-007                     level=54                         vth0=0.11074668 lvth0=-2.6843719e-008            wvth0=-4.761698e-008             pvth0=1.8250804e-014 k2=-0.0084341095              lk2=-1.8843098e-009            wk2=2.1328377e-009 pk2=1.325906e-015              u0=0.12739866                 lu0=-1.930754e-008 wu0=-3.4070993e-008            pu0=9.6141248e-015             ua=1.4796784e-009 lua=-3.4930866e-016            wua=-4.1931019e-016            pua=-1.1435405e-022 ub=5.7724877e-018             lub=-1.5031821e-024            wub=-2.0575499e-024 pub=9.5844332e-031             uc=-2.8013653e-011            luc=-8.0661223e-019 wuc=-1.0867519e-017            puc=9.1378723e-024             vsat=127200 a0=19.100336                  la0=-1.2926907e-005            wa0=-9.4919347e-006 pa0=8.1170767e-012             ags=6.5465836                  lags=-1.7197721e-006 wags=-1.7707972e-006            pags=7.0832168e-013             keta=-0.091894017 lketa=3.9120899e-008             wketa=-4.1480067e-009            pketa=1.9592862e-015 voff=-0.20769548                lvoff=2.8895946e-008             wvoff=6.6452575e-008 pvoff=-2.9359007e-014            minv=0.16393416                 lminv=-5.5069645e-007 wminv=-5.7337529e-007            pminv=5.0802247e-013             etab=-0.033219332 wetab=1.5003660e-008             cit=0.0018880935               lcit=1.3245229e-009 wcit=1.1665944e-009             pcit=-7.2649291e-016            pdiblc2=0.050933273 lpdiblc2=-6.7382531e-009            wpdiblc2=-9.3334002e-009            ppdiblc2=-1.0570193e-016 agidl=-7.4906262e-005            lagidl=3.1400577e-011             wagidl=7.3282006e-011 pagidl=-2.8614700e-017            aigbacc=0.015371067                laigbacc=-7.8653120e-010 waigbacc=-1.2421864e-009            paigbacc=7.1259727e-016             bigbacc=0.0058832969 lbigbacc=-3.8688404e-010            wbigbacc=-8.3244810e-010            pbigbacc=3.6461227e-016 aigc=0.011979899                laigc=2.3016208e-011             waigc=5.5659533e-011 paigc=-6.1943705e-017            bigc=0.0015455                  aigsd=0.010308138 laigsd=2.6688487e-011             waigsd=4.0474628e-011             paigsd=-1.3789945e-017 bigsd=0.00063047289              lbigsd=3.0452875e-011             wbigsd=3.7961803e-011 pbigsd=-1.6627270e-017            ute=-0.56051364                lute=-4.2169020e-007 wute=-3.3030799e-007            pute=2.4133294e-013             kt1=-0.20483914 lkt1=-5.663356e-008             wkt1=1.4422737e-008             pkt1=-5.0713172e-015 kt2=1.9442222e-006             lkt2=-7.2658773e-009            wkt2=-5.8111422e-009 pkt2=3.0261631e-015             ua1=6.5615174e-009             lua1=7.7471883e-018 wua1=-1.0977978e-015            pua1=-2.3254424e-022            ub1=-8.9589644e-019 lub1=-3.4406346e-024            wub1=-2.5974521e-024            pub1=2.5433784e-030 uc1=4.065248e-011              luc1=-2.2110487e-017            wuc1=-3.2843757e-017 puc1=7.4371401e-024             at=223608.12                  lat=-0.096004301 wat=-0.039305141               pat=3.7087125e-008             tvoff=8.1551389e-005 ltvoff=2.6838937e-010             wtvoff=3.2420744e-009             ptvoff=-1.4177716e-015 lvsat=0                          wvsat=0                          pvsat=0 vsat_mc=1907.74                    lvsat_mc=-0.00169407                wvsat_mc=-0.00481485 pvsat_mc=4.27558e-09 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na12_mac.6 nmos ( lmin=2.7e-07                    lmax=4.5e-007                   wmin=5.4e-007 wmax=9e-007                     level=54                         vth0=0.14636137 lvth0=-4.2442953e-008            wvth0=-8.7528933e-008            pvth0=3.5732239e-014 k2=-0.019349047               lk2=2.8964327e-009             wk2=7.7743921e-009 pk2=-1.1450949e-015            u0=0.10858568                 lu0=-1.1067455e-008 wu0=-2.8600105e-008            pu0=7.2178761e-015             ua=1.5479456e-009 lua=-3.7920967e-016            wua=-8.1179057e-016            pua=5.7552361e-023 ub=2.5873826e-018             lub=-1.0810611e-025            wub=-2.5318709e-025 pub=1.6813243e-031             uc=-1.545238e-010             luc=5.4604830e-017 wuc=8.5515373e-017             puc=-3.3077834e-023            vsat=174372.19 a0=-34.271222                 la0=1.0449836e-005             wa0=2.6194926e-005 pa0=-7.5137684e-012            ags=5.7797173                  lags=-1.3838847e-006 wags=-1.5055189e-006            pags=5.9212981e-013             keta=-0.079503573 lketa=3.3693885e-008             wketa=4.1168654e-008             pketa=-1.7889411e-014 voff=-0.20137308                lvoff=2.6126734e-008             wvoff=6.2802782e-008 pvoff=-2.7760398e-014            minv=-2.9154127                 lminv=7.9805748e-007 wminv=1.7619562e-006             pminv=-5.1485273e-013            etab=-0.11731572 wetab=7.5720742e-008             cit=0.0042878634               lcit=2.7342364e-010 wcit=2.5244874e-009             pcit=-1.32125e-015              pdiblc2=0.066916511 lpdiblc2=-1.3738911e-008            wpdiblc2=-2.3485613e-008            ppdiblc2=6.0929674e-015 agidl=-2.1702234e-005            lagidl=8.0972127e-012             wagidl=2.3326882e-011 pagidl=-6.7343551e-018            aigbacc=0.012157289                laigbacc=6.2110347e-010 waigbacc=1.4876923e-009             paigbacc=-4.8308959e-016            bigbacc=0.0011956944 lbigbacc=1.6662858e-009             wbigbacc=3.4467008e-009             pbigbacc=-1.5096550e-015 aigc=0.012263852                laigc=-1.0135500e-010            waigc=-1.9220645e-010 paigc=4.6621596e-017             bigc=0.0017135416               aigsd=0.010341972 laigsd=1.1869218e-011             waigsd=2.6781621e-011             paigsd=-7.7924076e-018 bigsd=0.0007                     ute=-2.2504678                 lute=3.1850973e-007 wute=4.3843317e-007             pute=-9.5375687e-014            kt1=-0.29492087 lkt1=-1.7177759e-008            wkt1=-1.2204436e-007            pkt1=5.4701269e-014 kt2=-0.024811809               lkt2=3.6025466e-009             wkt2=8.2315919e-009 pkt2=-3.1245544e-015            ua1=7.9085476e-009             lua1=-5.8225206e-016 wua1=-1.2858232e-015            pua1=-1.5018910e-022            ub1=-1.3498692e-017 lub1=2.0793897e-024             wub1=4.1115958e-024             pub1=-3.9518454e-031 uc1=1.0800995e-010             luc1=-5.161306e-017             wuc1=-1.4976339e-016 puc1=5.8647939e-023             at=-32537.089                 lat=0.0161873 wat=0.085330697                pat=-1.750337e-008             tvoff=0.00024637553 ltvoff=1.9619639e-010             wtvoff=-7.0516293e-010            ptvoff=3.1111832e-016 lvsat=-0.020661421               wvsat=-0.017233504               pvsat=7.5482748e-009 letab=3.6834219e-008             petab=-2.6594082e-014            lbigc=-7.3602226e-011 wbigc=-1.5224570e-010            pbigc=6.6683616e-017             vth0_mc=-0.00731002 lvth0_mc=3.20182e-09                wvth0_mc=1.18172e-08                pvth0_mc=-5.17594e-15 vsat_mc=-3359.84                   lvsat_mc=0.00061315                 wvsat_mc=0.0140067 pvsat_mc=-3.96824e-09 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na12_mac.7 nmos ( lmin=9e-007                     lmax=9.019e-06                  wmin=4.5e-07 wmax=5.4e-007                   level=54                         vth0=-0.022659328 lvth0=1.2079268e-007             wvth0=2.0726947e-008             pvth0=-5.8366442e-014 k2=0.0068808191               lk2=-2.0159896e-008            wk2=-2.8602543e-009 pk2=8.3128294e-015             u0=0.070303845                lu0=1.404664e-008 wu0=-4.6375602e-009            pu0=-7.0518394e-015            ua=4.6934416e-009 lua=-4.4105938e-015            wua=-1.7950275e-015            pua=1.766558e-021 ub=-4.0734115e-018            lub=7.3416212e-024             wub=2.705824e-024 pub=-3.3269308e-030            uc=-7.234262e-011             luc=-5.3145267e-017 wuc=1.5547620e-017             puc=3.5750945e-023             vsat=127200 a0=7.7523443                  la0=-8.2854168e-006            wa0=1.1771581e-006 pa0=1.6107197e-012             ags=0.78150836                 lags=3.0695067e-006 wags=1.848115e-007              pags=-8.4801981e-013            keta=-0.13401217 lketa=9.2760100e-008             wketa=4.1492611e-008             pketa=-4.7435682e-014 voff=-0.11212361                lvoff=-2.0922814e-008            wvoff=8.6692132e-009 pvoff=2.8158292e-015             minv=-0.3430738                 lminv=-1.8057689e-006 wminv=-6.2195147e-008            pminv=9.8518586e-013             etab=-0.16148994 wetab=8.5039413e-008             cit=0.0084541299               lcit=-4.4122381e-009 wcit=-2.3952208e-009            pcit=2.3851409e-015             pdiblc2=0.028111965 lpdiblc2=6.7113578e-009             wpdiblc2=-4.1044237e-009            ppdiblc2=-1.027655e-015 agidl=-1.1669768e-005            lagidl=1.8032308e-010             wagidl=8.4991874e-012 pagidl=-8.3059329e-017            aigbacc=0.012676439                laigbacc=5.1204099e-009 waigbacc=2.3289809e-010             paigbacc=-2.5159829e-015            bigbacc=0.0035461961 lbigbacc=6.9638179e-009             wbigbacc=2.4130098e-010             pbigbacc=-3.4692215e-015 aigc=0.012328789                laigc=-4.4470078e-010            waigc=-5.7077471e-011 paigc=1.2438169e-016             bigc=0.0015455                  aigsd=0.010482857 laigsd=-1.0757600e-010            waigsd=-3.6904528e-010            paigsd=3.3845967e-016 bigsd=0.00078281684              lbigsd=-7.3541352e-011            wbigsd=-2.9076003e-010 pbigsd=2.5819491e-016             ute=-1.2511939                 lute=2.9079682e-007 wute=-1.0937854e-007            pute=-8.9953885e-015            kt1=-0.0052487516 lkt1=2.3345595e-008             wkt1=-8.1171258e-008            pkt1=-6.0623467e-014 kt2=0.01193628                 lkt2=-2.0840899e-008            wkt2=-1.8794262e-008 pkt2=1.6180796e-014             ua1=1.14946e-008               lua1=-7.4894042e-015 wua1=-4.7269325e-015            pua1=4.6917766e-021             ub1=-2.3725519e-017 lub1=1.8983190e-023             wub1=1.0957562e-023             pub1=-1.0667986e-029 uc1=-1.9306654e-010            luc1=2.8131314e-017             wuc1=1.1348507e-016 puc1=-3.6616683e-023            at=-152036.41                 lat=0.15846811 wat=0.138305                   pat=-7.7442118e-008            tvoff=0.007417122 ltvoff=1.8503120e-009             wtvoff=4.1198950e-010             ptvoff=-3.3250227e-015 lvsat=0                          wvsat=0                          pvsat=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na12_mac.8 nmos ( lmin=4.5e-007                   lmax=9e-007                     wmin=4.5e-07 wmax=5.4e-007                   level=54                         vth0=0.14354388 lvth0=-2.6795764e-008            wvth0=-6.552425e-008             pvth0=1.822462e-014 k2=-0.021683628               lk2=5.2053326e-009             wk2=9.3670747e-009 pk2=-2.5450388e-015            u0=0.086857065                lu0=-6.5261922e-010 wu0=-1.1935282e-008            pu0=-5.7146211e-016            ua=-1.056028e-009 lua=6.9493518e-016             wua=9.6518553e-016             pua=-6.8451118e-022 ub=5.8477695e-018             lub=-1.4683875e-024            wub=-2.0986537e-024 pub=9.3944545e-031             uc=-2.4847155e-010            luc=1.0325722e-016 wuc=1.0950249e-016             puc=-4.7680981e-023            vsat=127200 a0=-17.201715                 la0=1.3873788e-005             wa0=1.0328985e-005 pa0=-6.5161027e-012            ags=6.801946                   lags=-2.2766419e-006 wags=-1.910225e-006             pags=1.0123726e-012             keta=-0.24770747 lketa=1.9372153e-007             wketa=8.0926141e-008             pketa=-8.2452657e-014 voff=-0.16635831                lvoff=2.7237604e-008             wvoff=4.3882481e-008 pvoff=-2.8453553e-014            minv=-5.1043186                 lminv=2.4222165e-006 wminv=2.3030907e-006             pminv=-1.1151880e-012            etab=-0.16148994 wetab=8.5039413e-008             cit=0.00066050747              lcit=2.5084986e-009 wcit=1.8368564e-009             pcit=-1.3729437e-015            pdiblc2=0.030782109 lpdiblc2=4.3402693e-009             wpdiblc2=1.6691351e-009             ppdiblc2=-6.1545752e-015 agidl=0.00033378773              lagidl=-1.2644318e-010            wagidl=-1.4986491e-010 pagidl=5.7567993e-017             aigbacc=0.021113493                laigbacc=-2.3716941e-009 waigbacc=-4.3775514e-009            paigbacc=1.5780962e-015             bigbacc=0.01662 lbigbacc=-4.6457200e-009            wbigbacc=-6.6946880e-009            pbigbacc=2.6899367e-015 aigc=0.011760342                laigc=6.0080036e-011             waigc=1.7553767e-010 paigc=-8.2180555e-017            bigc=0.0015455                  aigsd=0.010349374 laigsd=1.0956985e-011             waigsd=1.7959469e-011             paigsd=-5.2005443e-018 bigsd=0.0007                     ute=-1.0822111                 lute=1.4074011e-007 wute=-4.5461173e-008            pute=-6.5754008e-014            kt1=0.55958342 lkt1=-4.7822537e-007            wkt1=-4.0295198e-007            pkt1=2.2511781e-013 kt2=-0.028085707               lkt2=1.4698626e-008             wkt2=9.5247152e-009 pkt2=-8.9664557e-015            ua1=1.1978732e-009             lua1=1.6540895e-015 wua1=1.8307519e-015             pua1=-1.1314472e-021            ub1=-3.5199532e-018 lub1=1.0406470e-024             wub1=-1.1647171e-024            pub1=9.6598616e-032 uc1=-5.2574566e-011            luc1=-9.662556e-017             wuc1=1.8058211e-017 puc1=4.812237e-023              at=-193691.91                 lat=0.19545819 wat=0.18854067                 pat=-1.2205139e-007            tvoff=0.02272976 ltvoff=-1.1747310e-008            wtvoff=-9.1238472e-009            ptvoff=5.1428003e-015 lvsat=0                          wvsat=0                          pvsat=0 vsat_mc=-41924.7                   lvsat_mc=0.0372291                  wvsat_mc=0.0191177 pvsat_mc=-1.69765e-08 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na12_mac.9 nmos ( lmin=2.7e-07                    lmax=4.5e-007                   wmin=4.5e-07 wmax=5.4e-007                   level=54                         vth0=-0.064769824 lvth0=6.4445637e-008             wvth0=2.7748698e-008             pvth0=-2.2628931e-014 k2=-0.0026994677              lk2=-3.1097295e-009            wk2=-1.316278e-009 pk2=2.1342697e-015             u0=0.12380907                 lu0=-1.6837596e-008 wu0=-3.6912075e-008            pu0=1.0368373e-014             ua=4.1114261e-009 lua=-1.5684097e-015            wua=-2.2114509e-015            pua=7.0685559e-022 ub=6.8319978e-019             lub=7.9369406e-025             wub=7.8649674e-025 pub=-3.2425046e-031            uc=9.2520709e-011             luc=-4.6097387e-017 wuc=-4.9370926e-017            puc=2.1905576e-023             vsat=171131.67 a0=53.080433                  la0=-1.6909793e-005            wa0=-2.1499078e-005 pa0=7.4245888e-012             ags=0.019698                   lags=6.9398268e-007 wags=1.6394516e-006             pags=-5.4238575e-013            keta=0.029315748 lketa=7.2385357e-008             wketa=-1.8246695e-008            pketa=-3.9014955e-014 voff=0.084212911                lvoff=-8.2512591e-008            wvoff=-9.3127167e-008 pvoff=3.1556673e-014             minv=3.0840663                  lminv=-1.1642961e-006 wminv=-1.5137593e-006            pminv=5.5639233e-013             etab=0.0029595371 wetab=1.0050451e-008             cit=0.027133683                lcit=-9.0867521e-009 wcit=-9.9493299e-009            pcit=3.7894059e-015             pdiblc2=0.071621109 lpdiblc2=-1.3547212e-008            wpdiblc2=-2.6054324e-008            ppdiblc2=5.9882999e-015 agidl=0.00011023707              lagidl=-2.8527994e-011            wagidl=-4.8711979e-011 pagidl=1.3263008e-017             aigbacc=0.017905618                laigbacc=-9.6664459e-010 waigbacc=-1.6508953e-009            paigbacc=3.8382085e-016             bigbacc=0.019778111 lbigbacc=-6.0289727e-009            wbigbacc=-6.6992987e-009            pbigbacc=2.6919562e-015 aigc=0.010023414                laigc=8.2085461e-010             waigc=1.0310726e-009 paigc=-4.5690485e-016            bigc=-0.00047380867             aigsd=0.01189402 laigsd=-6.6559779e-010            waigsd=-8.2063670e-010            paigsd=3.6210458e-016 bigsd=0.0018793849               lbigsd=-5.1657058e-010            wbigsd=-6.4394415e-010 pbigsd=2.8204754e-016             ute=-0.96050413                lute=8.7432450e-008 wute=-2.6588700e-007            pute=3.0792505e-014             kt1=-1.377041 lkt1=3.7001611e-007             wkt1=4.6879322e-007             pkt1=-1.5670658e-013 kt2=0.035672847                lkt2=-1.3227620e-008            wkt2=-2.4793030e-008 pkt2=6.0647168e-015             ua1=1.38279e-008               lua1=-3.8778620e-015 wua1=-4.5177894e-015            pua1=1.6492139e-021             ub1=-9.5281198e-018 lub1=3.6722240e-024             wub1=1.9436634e-024             pub1=-1.2648721e-030 uc1=-9.5427344e-010            luc1=2.9831855e-016             wuc1=4.3024335e-016 puc1=-1.3241472e-022            at=418438.09                  lat=-0.072654747 wat=-0.16090176                pat=3.1004388e-008             tvoff=-0.015306135 ltvoff=4.9124115e-009             wtvoff=7.7865077e-009             ptvoff=-2.2639351e-015 lvsat=-0.01924207                wvsat=-0.015464176               pvsat=6.7733091e-009 letab=-7.2028871e-008            petab=3.2845165e-014             lbigc=8.8445720e-010 wbigc=1.0420476e-009             pbigc=-4.5641683e-016            vth0_mc=0.0869559 lvth0_mc=-3.80865e-08               wvth0_mc=-3.96518e-08               pvth0_mc=1.73675e-14 vsat_mc=135246                     uc1_ff=-0                         luc1_ff=0 wuc1_ff=0                          puc1_ff=0.35e-23                   lvsat_mc=-0.0403717 wvsat_mc=-0.0616723                 pvsat_mc=1.84095e-08 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_na18_mac.global nmos ( modelid=15                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=0                          igbmod=0 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_na18'            permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=3.36e-009                  toxm=3.36e-009                  dtox=1.9844e-010 epsrox=3.9                        wint=0                          lint=0 ll=0                          wl=0                          lln=1 wln=1                          lw=0                          ww=0 lwn=1                          wwn=1                          lwl=0 wwl=0                          llc=0                          wlc=0 lwc=0                          wwc=0                          lwlc=0 wwlc=0                          xl=1e-008                     xw=0 dlc=3.542614e-008              dwc=0                          xpart=1 toxref=3e-009                     dlcig=2.5e-009                   k1=0.054 k3=-8.2825                    k3b=-4.2795                    w0=0 dvt0=0.0050825                  dvt1=45.501                     dvt2=0.185 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.062479                   voffl=-5e-009                    dvtp0=0 dvtp1=4                          lpe0=-4.24e-007                 lpeb=-1e-007 xj=6.7e-008                   ngate=3e+021                     ndep=1e+017 nsd=1e+020                     phin=0.19                       cdsc=0 cdscb=0                          cdscd=0                          nfactor=0.53 ud=0                          lud=0                          wud=0 pud=0                          a1=0                          a2=1 b0=0                          b1=0                          dwg=0 dwb=0                          pdiblc1=0                          pdiblcb=0 drout=0.56                       pvag=0.3                        delta=0.01 pscbe1=9.264e+008                 pscbe2=1e-020                     fprout=100 pdits=0                          pditsd=0                          pditsl=0 rsh=18.0                       rdsw=217.15                     prwg=0 prwb=0                          wr=1                          alpha0=0 alpha1=0.00035                    beta0=7                          agidl=1.4314e-011 bgidl=2.3e+009                   cgidl=0.5                        egidl=0.8 aigbacc=0.01238                    bigbacc=0.006109                   cigbacc=0.2809 nigbacc=4.05                       aigbinv=0.0111                     bigbinv=0.000949 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1 aigc=0.009898                   bigc=0.001383                   cigc=1.515e-005 aigsd=0.0086                     bigsd=0.0004353                  cigsd=3.925e-020 nigc=1                          poxedge=1                          pigcd=1.672 ntox=1                          xrcrg1=12                         xrcrg2=1 vfbsdoff=0                          lvfbsdoff=0                          wvfbsdoff=0 pvfbsdoff=0                          cgso=4.925043e-011              cgdo=4.925043e-011 cgbo=0                          cgdl=3.247859e-010              cgsl=3.247859e-010 clc=0                          cle=0.6                        cf='8.050e-11+7.81e-11*ccoflag_na18' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=16.193                     noff=3.9                        voffcv=-0.004675 kt1l=0                          prt=0                          fnoimod=1.000000e+00 tnoimod=0                          em=1.300000e+06               ef=1.050000e+00 noia=0                          noib=0                          noic=0 lintnoi=-1.000000e-07              jss=1.60e-06                   jsd=1.60e-06 jsws=1.57e-12                   jswd=1.57e-12                   jswgs=1.57e-12 jswgd=1.57e-12                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=19.65                      bvd=19.65 xjbvs=1                          xjbvd=1                          jtsswgs=1.6e-010 jtsswgd=1.6e-010                   njtsswg=20                         xtsswgs=0.69066 xtsswgd=0.69066                    tnjtsswg=1                          vtsswgs=10 vtsswgd=10                         pbs=0.512                      pbd=0.512 cjs=0.000161                   cjd=0.000161                   mjs=0.292 mjd=0.292                      pbsws=0.3                        pbswd=0.3 cjsws=2.08e-010                  cjswd=2.08e-010                  mjsws=0.039 mjswd=0.039                      pbswgs=0.791                      pbswgd=0.791 cjswgs=1.62e-010                  cjswgd=1.62e-010                  mjswgs=0.385 mjswgd=0.385                      tpb=0.0014                     tcj=0.0012 tpbsw=0.0013                     tcjsw=0.00034                    tpbswg=0.0022 tcjswg=0.0015                     xtis=3                          xtid=3 dmcg=6.7e-008                   dmci=6.7e-008                   dmdg=0 dmcgt=0                          dwj=0                          xgw=0 xgl=2.64e-09                   rshg=16.42                      gbmin=1e-012 rbpb=50                         rbpd=50                         rbps=50 rbdb=50                         rbsb=50                         ngcon=1 lnfactor=0                          pnfactor=0                          rdw=0 rsw=0                          wnfactor=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.7 sigma_factor='sigma_factor_na18' ccoflag='ccoflag_na18' rcoflag='rcoflag_na18' rgflag='rgflag_na18' mismatchflag='mismatchflag_mos_na18' globalflag='globalflag_mos_na18' totalflag='totalflag_mos_na18' global_factor='global_factor_na18' local_factor='local_factor_na18' sigma_factor_flicker='sigma_factor_flicker_na18' noiseflag='noiseflagn_na18' noiseflag_mc='noiseflagn_na18_mc' delvto=0 mulu0=1 dlc_fmt=2 par1_io='par1_io' par2_io='par2_io' par3_io='par3_io' par4_io='par4_io' par5_io='par5_io' par6_io='par6_io' par7_io='par7_io' par8_io='par8_io' par9_io='par9_io' par10_io='par10_io' par11_io='par11_io' par12_io='par12_io' par13_io='par13_io' par14_io='par14_io' par15_io='par15_io' par16_io='par16_io' par17_io='par17_io' par18_io='par18_io' par19_io='par19_io' par20_io='par20_io' w1_io='2.0857*0.40825' w2_io='0.67082*-0.40825' w3_io='0.54772*0.26807' w4_io='0.54772*-0.6902' w5_io='0.54772*-0.32981' w6_io='0.54772*0.098267' tox_c='toxn_na18'                dxl_c='dxln_na18'                dxw_c='dxwn_na18' cj_c='cjn_na18'                 cjsw_c='cjswn_na18'               cjswg_c='cjswgn_na18' cgo_c='cgon_na18'                cgl_c='cgln_na18'                ddlc_c='ddlcn_na18' dvth_c='dvthn_na18'               dlvth_c='dlvthn_na18'              dwvth_c='dwvthn_na18' dpvth_c='dpvthn_na18'              cf_c='cfn_na18'                 du0_c='du0n_na18' dlu0_c='dlu0n_na18'               dwu0_c='dwu0n_na18'               dpu0_c='dpu0n_na18' dvsat_c='dvsatn_na18'              dlvsat_c='dlvsatn_na18'             dwvsat_c='dwvsatn_na18' dpvsat_c='dpvsatn_na18'             dk2_c='dk2n_na18'                drdsw_c='drdswn_na18' dvoff_c='dvoffn_na18'              dlvoff_c='dlvoffn_na18'             dwvoff_c='dwvoffn_na18' dpvoff_c='dpvoffn_na18'             dpdiblc2_c='dpdiblc2n_na18'           dlpdiblc2_c='dlpdiblc2n_na18' dwpdiblc2_c='dwpdiblc2n_na18'          dppdiblc2_c='dppdiblc2n_na18'          dags_c='dagsn_na18' dlags_c='dlagsn_na18'              dwags_c='dwagsn_na18'              dpags_c='dpagsn_na18' dnfactor_c='dnfactorn_na18'           dlnfactor_c='dlnfactorn_na18'          dwnfactor_c='dwnfactorn_na18' dpnfactor_c='dpnfactorn_na18'          dcit_c='dcitn_na18'               dlcit_c='dlcitn_na18' dwcit_c='dwcitn_na18'              dpcit_c='dpcitn_na18'              deta0_c='deta0n_na18' dleta0_c='dleta0n_na18'             dweta0_c='dweta0n_na18'             dpeta0_c='dpeta0n_na18' dub1_c='dub1n_na18'               dlk2_c='dlk2n_na18'               dwk2_c='dwk2n_na18' dpk2_c='dpk2n_na18'               dkt1_c='dkt1n_na18'               dlkt2_c='dlkt2n_na18' dla0_c='dla0n_na18'               dwa0_c='dwa0n_na18'               dluc_c='dlucn_na18' dlketa_c='dlketan_na18'             monte_flag_c='monte_flagn_na18'        c1f_c='c1fn_na18' c2f_c='c2fn_na18'                c3f_c='c3fn_na18' global_mc='global_mc_flag_na18' tox_g='toxn_na18_ms_global'      dxl_g='dxln_na18_ms_global'      dxw_g='dxwn_na18_ms_global' cj_g='cjn_na18_ms_global'       cjsw_g='cjswn_na18_ms_global' cjswg_g='cjswgn_na18_ms_global'    cgo_g='cgon_na18_ms_global'      cgl_g='cgln_na18_ms_global' dvth_g='dvthn_na18_ms_global'     dlvth_g='dlvthn_na18_ms_global' dwvth_g='dwvthn_na18_ms_global'    dpvth_g='dpvthn_na18_ms_global' cf_g='cfn_na18_ms_global'       du0_g='du0n_na18_ms_global' dlu0_g='dlu0n_na18_ms_global'     dwu0_g='dwu0n_na18_ms_global' dpu0_g='dpu0n_na18_ms_global'     dvsat_g='dvsatn_na18_ms_global' dlvsat_g='dlvsatn_na18_ms_global'   dwvsat_g='dwvsatn_na18_ms_global' dpvsat_g='dpvsatn_na18_ms_global'   dk2_g='dk2n_na18_ms_global' dlvoff_g='dlvoffn_na18_ms_global'   dppdiblc2_g='dppdiblc2n_na18_ms_global' dags_g='dagsn_na18_ms_global'     dwags_g='dwagsn_na18_ms_global' deta0_g='deta0n_na18_ms_global'    dlk2_g='dlk2n_na18_ms_global' dwk2_g='dwk2n_na18_ms_global'     dpk2_g='dpk2n_na18_ms_global' dkt1_g='dkt1n_na18_ms_global'     dlkt2_g='dlkt2n_na18_ms_global' dla0_g='dla0n_na18_ms_global'     dwa0_g='dwa0n_na18_ms_global' dluc_g='dlucn_na18_ms_global'     dlketa_g='dlketan_na18_ms_global' monte_flag_g='monte_flagn_na18_ms_global'                                      ddlc_g='ddlcn_na18_ms_global' weight1=-3.1983125 weight2=1.5975625 weight3=-1.038375 weight4=-0.625 weight5=-0.4297125 tox_1=1.2526e-011 tox_2=-2.6961e-011 tox_3=-1.0998e-012 tox_4=9.4257e-011 tox_5=4.0716e-012 dxl_1=7.5174e-010 dxl_2=-1.618e-009 dxl_3=-6.6005e-011 dxl_4=-5.6569e-009 dxl_5=2.4436e-010 dxw_1=-1.2161e-009 dxw_2=-2.3698e-009 dxw_3=-1.3015e-009 dxw_4=-2.1115e-024 dxw_5=-1.1627e-008 cj_1=1.0896e-006 cj_2=-1.1204e-007 cj_3=4.5396e-007 cj_4=2.0024e-021 cj_5=-1.431e-007 cjsw_1=1.4077e-012 cjsw_2=-1.4475e-013 cjsw_3=5.8648e-013 cjsw_4=-2.9972e-028 cjsw_5=-1.8487e-013 cjswg_1=1.0964e-012 cjswg_2=-1.1274e-013 cjswg_3=4.5678e-013 cjswg_4=5.2561e-028 cjswg_5=-1.4399e-013 cgo_1=-3.3333e-013 cgo_2=3.4274e-014 cgo_3=-1.3887e-013 cgo_4=4.3203e-028 cgo_5=4.3775e-014 cgl_1=-2.1982e-012 cgl_2=2.2602e-013 cgl_3=-9.1577e-013 cgl_4=3.2719e-027 cgl_5=2.8868e-013 dvth_1=0.006065 dvth_2=0.0034522 dvth_3=0.0032314 dvth_4=-3.8046e-018 dvth_5=-0.0016707 dlvth_1=1.3793e-009 dlvth_2=8.4963e-010 dlvth_3=5.4735e-010 dlvth_4=1.1923e-025 dlvth_5=-3.7158e-010 dwvth_1=3.7255e-010 dwvth_2=1.5998e-010 dwvth_3=1.4975e-010 dwvth_4=4.9101e-025 dwvth_5=-8.7014e-011 dpvth_1=4.8676e-017 dpvth_2=2.0468e-016 dpvth_3=-9.0892e-017 dpvth_4=-9.9193e-033 dpvth_5=-3.4886e-017 cf_1=-5.4482e-013 cf_2=5.6021e-014 cf_3=-2.2698e-013 cf_4=1.0968e-027 cf_5=7.155e-014 du0_1=4.8192e-005 du0_2=0.00047724 du0_3=0.00013197 du0_4=-1.5639e-019 du0_5=-0.00011294 dlu0_1=-1.7706e-011 dlu0_2=1.1738e-010 dlu0_3=2.1062e-011 dlu0_4=5.9835e-027 dlu0_5=-2.3406e-011 dwu0_1=3.0143e-013 dwu0_2=7.9941e-011 dwu0_3=1.5712e-013 dwu0_4=-1.9145e-026 dwu0_5=-1.8178e-011 dpu0_1=-1.2201e-017 dpu0_2=1.0069e-016 dpu0_3=-2.1616e-018 dpu0_4=3.3721e-032 dpu0_5=-2.0657e-017 dvsat_1=-966.86 dvsat_2=99.417 dvsat_3=-402.8 dvsat_4=-1.7393e-012 dvsat_5=126.97 dlvsat_1=0.00054684 dlvsat_2=-7.7595e-005 dlvsat_3=0.00042603 dlvsat_4=-5.1274e-019 dlvsat_5=-8.9805e-005 dwvsat_1=-0.00024778 dwvsat_2=1.1234e-005 dwvsat_3=2.8912e-005 dwvsat_4=-5.4722e-020 dwvsat_5=2.0547e-005 dpvsat_1=1.0777e-010 dpvsat_2=4.7294e-012 dpvsat_3=-1.0178e-010 dpvsat_4=1.3419e-025 dpvsat_5=-8.4078e-013 dk2_1=0.00013668 dk2_2=-1.7758e-005 dk2_3=9.13e-005 dk2_4=3.0668e-020 dk2_5=-2.1068e-005 dlvoff_1=-2.1765e-010 dlvoff_2=-3.4598e-011 dlvoff_3=4.3789e-010 dlvoff_4=2.7605e-025 dlvoff_5=-1.9391e-011 dppdiblc2_1=4.2274e-018 dppdiblc2_2=-1.8591e-018 dppdiblc2_3=1.4975e-017 dppdiblc2_4=-7.1959e-033 dppdiblc2_5=-1.7545e-018 dags_1=-0.002906 dags_2=0.00062643 dags_3=-0.0042499 dags_4=-3.596e-018 dags_5=0.00065749 dwags_1=1.39e-009 dwags_2=-5.7462e-011 dwags_3=-2.1375e-010 dwags_4=-1.0871e-024 dwags_5=-1.1059e-010 deta0_1=-0.0004502 deta0_2=4.4867e-005 deta0_3=-0.00017434 deta0_4=2.7218e-019 deta0_5=5.7923e-005 dlk2_1=4.5329e-011 dlk2_2=-3.8768e-013 dlk2_3=-2.0758e-011 dlk2_4=-5.0997e-026 dlk2_5=-2.3549e-012 dwk2_1=4.2316e-011 dwk2_2=4.1955e-012 dwk2_3=-6.1655e-011 dwk2_4=1.5331e-026 dwk2_5=1.6389e-012 dpk2_1=1.4503e-016 dpk2_2=-1.4913e-017 dpk2_3=6.042e-017 dpk2_4=1.3354e-031 dpk2_5=-1.9046e-017 dkt1_1=-0.0022058 dkt1_2=0.00015559 dkt1_3=-0.00025824 dkt1_4=1.1147e-018 dkt1_5=0.00022971 dlkt2_1=1.6324e-011 dlkt2_2=2.5948e-012 dlkt2_3=-3.2842e-011 dlkt2_4=7.5187e-027 dlkt2_5=1.4543e-012 dla0_1=7.8562e-008 dla0_2=-5.2293e-009 dla0_3=6.3016e-009 dla0_4=1.6764e-022 dla0_5=-7.9187e-009 dwa0_1=-1.783e-008 dwa0_2=-3.0324e-010 dwa0_3=1.2393e-008 dwa0_4=3.754e-023 dwa0_5=5.4259e-010 dluc_1=5.4412e-019 dluc_2=8.6494e-020 dluc_3=-1.0947e-018 dluc_4=7.0457e-034 dluc_5=4.8477e-020 dlketa_1=-2.7206e-010 dlketa_2=-4.3247e-011 dlketa_3=5.4736e-010 dlketa_4=2.4041e-026 dlketa_5=-2.4239e-011 monte_flag_1=0.0939675 monte_flag_2=-0.20225 monte_flag_3=-0.00825062 monte_flag_4=-0.707113 monte_flag_5=0.030545 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.999982526 b_4=-4.20e-05                  c_4=-1.11e-04                  d_4=-1.04e-03 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=5.0e-06                    g_4_2=1.04988e-08 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.00185                    mis_a_2=-0.015                     mis_a_3=-0.035 mis_b_1=0.0010                     mis_b_2=0.16                       mis_b_3=0.01 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.002                      mis_d_2=0                          mis_d_3=0 mis_e_1=0.0017                     mis_e_2=0                          mis_e_3=0.23 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=0                          xl0=1e-8 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0                       bidirectionflag=1 designflag=1 cf0=8.050e-11                  cco=7.81e-11 noimod=1                          noic2='2.236'                    noic3='0.8' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.533e-6             sbref0=0.533e-6 samax=10e-6               sbmax=10e-6 samin=0.135e-6            sbmin=0.135e-6 rllodflag=0                   lreflod=1e-6                llodref=0.1 lod_clamp=-1e90 wlod0=1e-8 ku00=-3.0e-8             lku00=4e-6             wku00=0e-6 pku00=0.04e-11            tku00=0.8              llodku00=1 wlodku00=1                   kvsat0=0 kvth00=18.5e-9             lkvth00=14.0e-7          wkvth00=1.5e-6 pkvth00=0e-13               llodvth0=1                wlodvth0=1 stk20=7.5e-10             lodk20=1                steta00=-1.4e-9 lodeta00=1 wlod00=0 ku000=0e-8               lku000=0e-6               wku000=0e-6       		pku000=0.00e-11 llodku000=1                  wlodku000=1 kvth000=0e-8               lkvth000=-0e-15             wkvth000=-0e-15     		pkvth000=0 llodvth00=1                  wlodvth00=1                  steta000=-0e-9 stk200=0                  lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=0                wku01=0 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=0                wkvth01=0 pkvth01=0                   llodvth1=1                wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=0                   lku02=0                wku02=0 pku02=0                   tku02=0                llodku02=1 wlodku02=1                   kvsat2=1 kvth02=0                   lkvth02=0                wkvth02=0 pkvth02=0                   llodvth2=1                wlodvth2=1 stk22=0                   lodk22=1                steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0                pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0                   lku03=0                wku03=0 pku03=0                   tku03=0                llodku03=1 wlodku03=1                   kvsat3=0 kvth03=0                   lkvth03=0                wkvth03=0 pkvth03=0                   llodvth3=1                wlodvth3=1 stk23=0                   lodk23=1                steta03=0 lodeta03=1 wlod03=0 ku003=0.0e-2              lku003=-0.0e-8              wku003=0         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=5.33e-7             sa_b1=1.35e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.98e-7             spamax=1.6e-6              spamin=1.98e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=0.05                wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl=1.5e-6              ldplkvth0=0.8                 pkvth0dpl=0.0e-19 ku0dpl=0.20                wku0dpl=-3e-8               wdplku0=1 lku0dpl=6e-6                ldplku0=0.8                 pku0dpl=0.0e-11 keta0dpl=0                   wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=0                  wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx=0                   wku0dpx=0e-9                wdpxku0=1 lku0dpx=0e-8                ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=0                   wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps=0                   wku0dps=-0.0e-9             wdpsku0=1 lku0dps=0e-15               ldpsku0=2.0                 pku0dps=0e-23 keta0dps=0                   wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=-0.007              wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa=-1e-8               ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa=-0.02               wku0dpa=2e-9                wdpaku0=1 lku0dpa=-4.0e-8             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0.0                 wka0dpa=0                   wdpaka0=1 lka0dpa=0.0e-7              ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                   wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.31e-7             spbmax='1.6e-6+1.2e-6+0.2e-6'    spbmin='1.98e-7+1.98e-7+0.2e-6' pse_mode=1 kvth0dp2=0                   wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0e-9                ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.0                 wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=0e-5                ldp2ku0=0.5                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0                   wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1e-6 kvth0enx=0           	 wkvth0enx=0                   wenxkvth0=1 lkvth0enx=0          	 lenxkvth0=1                   pkvth0enx=0 ku0enx=0         		 wku0enx=0      		 wenxku0=1 lku0enx=0          	 lenxku0=1                   pku0enx=0 keta0enx=0                   wketa0enx=0                   wenxketa0=1 ka0enx=0                   wka0enx=0                   wenxka0=1 lka0enx=0          	 lenxka0=1                   pka0enx=0 kvsatenx=0                   wenx=0                   ku0enx0=0 eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0          	 wkvth0eny=0       		 wenykvth0=1 lkvth0eny=0        		 lenykvth0=1                   pkvth0eny=0 ku0eny=0          	 wku0eny=0        		 wenyku0=1 ku0eny0=0          	 wku0eny0=0                   weny0ku0=1 lku0eny=0       		 lenyku0=1                 	 pku0eny=0 keta0eny=0               	 wketa0eny=0                   wenyketa0=1 ka0eny=0              	 wka0eny=0             	 wenyka0=1 lka0eny=0      		 lenyka0=1                	 pka0eny=0 kvsateny=0               	 weny=0 kvth0eny1=0             	 wkvth0eny1=0        		 weny1kvth0=1 lkvth0eny1=0             	 leny1kvth0=1                  pkvth0eny1=0 ku0eny1=0        		 wku0eny1=0            	 weny1ku0=1 lku0eny1=0      		 leny1ku0=1                	 pku0eny1=0 keta0eny1=0              	 wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1                	 pka0eny1=0 kvsateny1=0               	 weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.8126e-5           ringxmin=0 kvth0rx=0              	 wkvth0rx=0          	 wrxkvth0=1 lkvth0rx=0              	 lrxkvth0=1                	 pkvth0rx=0 ku0rx=0              	 wku0rx=0           	 wrxku0=1 lku0rx=0        		 lrxku0=1                   pku0rx=0 keta0rx=0                	 wketa0rx=0                   wrxketa0=1 kvsatrx=0                	 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=1.6027e-5           ringymin=0 kvth0ry=0           	 wkvth0ry=0           	 wrykvth0=1 lkvth0ry=0              	 lrykvth0=1                 	 pkvth0ry=0 ku0ry=0          	 wku0ry=0           	 wryku0=1 lku0ry=0        		 lryku0=1                 	 pku0ry=0 keta0ry=0                	 wketa0ry=0                   wryketa0=1 kvsatry=0                   wry=0 kvth0ry0=0                	 ku0ry0=0 sfxref=8.26e-7           sfxmax=3e-6               minwodx=0.53e-6 sfxmin=0.189e-6 lrefodx=5e-8              lodxref=1                 wodx=1e-6 kvth0odxa=-0.200            lkvth0odxa=1.0e-13           lodxakvth0=2.0 wkvth0odxa=5.0e-12           wodxakvth0=2.0               pkvth0odxa=0.0e-16 ku0odxa=-1.20             lku0odxa=2.0e-13           lodxaku0=2.0 wku0odxa=5.0e-12           wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.0               wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0005           lkvth0odx1b=0.0e-7            lodx1bkvth0=0.5 wkvth0odx1b=-2.0e-15          wodx1bkvth0=2.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.00             lku0odx1b=0.0e-7            lodx1bku0=0.5 wku0odx1b=-1.5e-14          wodx1bku0=2.0               pku0odx1b=0.0e-16 sfyref=7.9e-7 sfymin=0.15e-6 sfymax=3e-6              minwody=0e-7              wody=1e-6 kvth0odya=-0.000            lkvth0odya=1.0e-13           lodyakvth0=2.0 wkvth0odya=0.0e-6            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=-2.00             lku0odya=2.0e-13           lodyaku0=2.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=0.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.00             lkvth0odyb=-3.0e-9           lodybkvth0=1.0 wkvth0odyb=-7.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=0.10              lku0odyb=0.0e-9            lodybku0=0.8 wku0odyb=-0.0e-5           wodybku0=1.0               pku0odyb=0.0e-13 web_mac=-0  wec_mac=-0 kvsatwe=-0 lodflag=1    pseflag=1 ceslflag=0 oseflag=1 wpeflag=0 )
.model nch_na18_mac.1 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-006                     wmax=0.00090001                 vth0=-0.1312 k2=0.0147                     minv=-0.21803                   cit=0.0001 voff=-0.118                     eta0=0.12                       etab=0.01 u0=0.042179                   ua=-3e-011                    ub=2.78e-018 uc=6.5485e-011                vsat=80000                      a0=6.7 ags=1.15                       keta=-0.028                     pclm=1 pdiblc2=0.0021                     tvoff=0.001824                   ltvoff=0 wtvoff=0                          ptvoff=0                          kt1=-0.17 kt2=-0.0024                    ute=-1.86                      ua1=8e-010 ub1=-2.6182e-018               uc1=-7.1e-011                  at=80000 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=0                          wk2=0 wvoff=0                          weta0=0                          wu0=0 wa0=0                          wags=0                          wpdiblc2=0 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wvsat=0                          pvsat=0 wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18_mac.2 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.13125028 k2=0.016409444                minv=-0.21803                   cit=0.0001 voff=-0.122525                  eta0=0.11698333                 etab=0.01 u0=0.041860993                ua=-3.2513889e-011            ub=2.7875417e-018 uc=7.2587842e-011             vsat=80000                      a0=7.0066944 ags=1.0557292                  keta=-0.024983333               pclm=0.84916667 pdiblc2=0.0013709722               tvoff=0.00145446                 ltvoff=3.32957e-009 wtvoff=0                          ptvoff=0                          kt1=-0.16874306 kt2=0.000274275                ute=-1.858014                  ua1=7.8464014e-010 ub1=-2.3012388e-018            uc1=-7.5005429e-011            at=80502.778 lvth0=4.5300278e-010             lk2=-1.5402094e-008            lvoff=4.077025e-008 leta0=2.7180167e-008             lu0=2.8652426e-009             lua=2.2650139e-017 lub=-6.7950417e-026            luc=-6.3996608e-017            la0=-2.7633169e-006 lags=8.4938021e-007             lketa=-2.7180167e-008            lpclm=1.3590083e-006 lpdiblc2=6.5685403e-009             lkt1=-1.1325069e-008            lkt2=-2.4095218e-008 lute=-1.789361e-008             lua1=1.3839235e-016             lub1=-2.8558201e-024 luc1=3.6088919e-017             lat=-0.0045300278              lvsat=0 lcit=0                          wvth0=0                          wk2=0 wvoff=0                          weta0=0                          wu0=0 wa0=0                          wags=0                          wpdiblc2=0 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wvsat=0                          pvsat=0 wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18_mac.3 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.13069722 k2=0.0060833333               minv=-0.21803                   cit=0.0001 voff=-0.1                       eta0=0.19558333                 etab=0.0061865139 u0=0.043737694                ua=-4.8611111e-012            ub=2.9392361e-018 uc=4.3058467e-011             vsat=78788.889                  a0=6.0552778 ags=1.7142361                  keta=-0.018805556               pclm=1.7513889 pdiblc2=0.0072708333               tvoff=0.00142102                 ltvoff=3.3901e-009 wtvoff=0                          ptvoff=0                          kt1=-0.18256944 kt2=-0.025206639               ute=-2.034125                  ua1=5.0579028e-010 ub1=-4.0326089e-018            uc1=-2.5047216e-011            at=149092.22 lvth0=-5.4802778e-010            lk2=3.2881667e-009             lvoff=0 leta0=-1.1508583e-007            lu0=-5.3158694e-010            lua=-2.7401389e-017 lub=-3.4251736e-025            luc=-1.0548439e-017            la0=-1.0412528e-006 lags=-3.4251736e-007            lketa=-3.8361944e-008            lpclm=-2.7401389e-007 lpdiblc2=-4.1102083e-009            lkt1=1.3700694e-008             lkt2=2.2025236e-008 lute=3.0086725e-007             lua1=6.431106e-016              lub1=2.7795969e-025 luc1=-5.4335447e-017            lat=-0.12867692                letab=6.9024099e-009 lvsat=0.0021921111               lcit=0                          wvth0=0 wk2=0                          wvoff=0                          weta0=0 wu0=0                          wa0=0                          wags=0 wpdiblc2=0                          pvth0=0                          pk2=0 pvoff=0                          peta0=0                          pu0=0 pags=0                          ppdiblc2=0                          wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18_mac.4 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.13870278 k2=0.012547222                minv=-0.51426806                cit=-0.0012789294 voff=-0.089861111               eta0=0.15083333                 etab=0.017626972 u0=0.041222222                ua=-3e-011                    ub=2.8277778e-018 uc=4.6510861e-011             vsat=81083.889                  a0=4.8972222 ags=1.9069444                  keta=-0.082388889               pclm=1.9055556 pdiblc2=0.0075555556               tvoff=-0.000205283               ltvoff=5.16277e-009 wtvoff=0                          ptvoff=0                          kt1=-0.18778361 kt2=0.01633425                 ute=-1.7603306                 ua1=1.5728347e-009 ub1=-5.3544e-018               uc1=-2.0737209e-010            at=83202.758 lvth0=8.1780278e-009             lk2=-3.7574722e-009            lvoff=-1.1051389e-008 leta0=-6.6308333e-008            lu0=2.2102778e-009             lub=-2.2102778e-025 luc=-1.4311549e-017            la0=2.2102778e-007             lags=-5.5256944e-007 lketa=3.0943889e-008             lpclm=-4.4205556e-007            lpdiblc2=-4.4205556e-009 lkt1=1.9384136e-008             lkt2=-2.3254333e-008            lute=2.4313056e-009 lua1=-5.1996785e-016            lub1=1.718712e-024              luc1=1.4439866e-016 lat=-0.056857407               letab=-5.5676897e-009            lvsat=-0.00030943889 lminv=3.2289948e-007             lcit=1.5030331e-009             wvth0=0 wk2=0                          wvoff=0                          weta0=0 wu0=0                          wa0=0                          wags=0 wpdiblc2=0                          pvth0=0                          pk2=0 pvoff=0                          peta0=0                          pu0=0 pags=0                          ppdiblc2=0                          wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18_mac.5 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.131375 k2=0.016125                   minv=-0.1725375                 cit=0.0001 voff=-0.123                     eta0=0.13312675                 etab=0.01 u0=0.04247375                 ua=-3.8e-011                  ub=2.8375e-018 uc=7.152075e-011              vsat=80000                      a0=7.0225 ags=1.1325                     keta=-0.031875                  pclm=1 pdiblc2=0.002125                   tvoff=0.00123                    ltvoff=0 wtvoff=5.346e-009                 ptvoff=0                          kt1=-0.17125 kt2=0.00088025                 ute=-1.865                     ua1=7.6451e-010 ub1=-2.50685e-018              uc1=-8.20675e-011              at=82500 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=1.575e-009                 wk2=-1.2825e-008 wminv=-4.094325e-007             wvoff=4.5e-008                   weta0=-1.1814075e-007 wu0=-2.65275e-009              wua=7.2e-017                   wub=-5.175e-025 wuc=-5.432175e-017             wa0=-2.9025e-006               wags=1.575e-007 wketa=3.4875e-008                wpdiblc2=-2.25e-010                 wkt1=1.125e-008 wkt2=-2.952225e-008             wute=4.5e-008                   wua1=3.1941e-016 wub1=-1.00215e-024              wuc1=9.96075e-017               wat=-0.0225 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wvsat=0                          pvsat=0 wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.6 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.13102934 k2=0.018431493                minv=-0.17283225                cit=0.0001 voff=-0.12909618                eta0=0.13099441                 etab=0.01 u0=0.042246432                ua=-3.9382639e-011            ub=2.8506979e-018 uc=8.090697e-011              vsat=80000                      a0=7.2999705 ags=1.0385434                  keta=-0.030460937               pclm=0.84288194 pdiblc2=0.0015279514               tvoff=0.00072232                 ltvoff=4.5742e-009 wtvoff=6.58924e-009               ptvoff=-1.12016e-014              kt1=-0.16999306 kt2=0.0047345602               ute=-1.8608018                 ua1=7.3182065e-010 ub1=-2.1329907e-018            uc1=-9.0283299e-011            at=83243.734 lvth0=-3.1143941e-009            lk2=-2.0781502e-008            lvoff=5.4926587e-008 leta0=1.9212414e-008             lu0=2.0481388e-009             lua=1.2457576e-017 lub=-1.1891323e-025            luc=-8.4569843e-017            la0=-2.5000091e-006 lags=8.4654894e-007             lketa=-1.2740703e-008            lpclm=1.4156337e-006 lpdiblc2=5.379408e-009              lkt1=-1.1325069e-008            lkt2=-3.4727335e-008 lute=-3.7825732e-008            lua1=2.9453108e-016             lub1=-3.368472e-024 luc1=7.4024346e-017             lat=-0.0067010436              lvsat=0 lminv=2.6557288e-009             lcit=0                          wvth0=-1.9884375e-009 wk2=-1.8198438e-008            wminv=-4.0677972e-007            wvoff=5.9140625e-008 weta0=-1.2609966e-007            wu0=-3.4689469e-009            wua=6.181875e-017 wub=-5.6840625e-025            wuc=-7.4872151e-017            wa0=-2.6394844e-006 wags=1.5467187e-007             wketa=4.9298438e-008             wpdiblc2=-1.4128125e-009 wkt1=1.125e-008                 wkt2=-4.0142566e-008            wute=2.509e-008 wua1=4.7537544e-016             wub1=-1.5142329e-024            wuc1=1.3750082e-016 wat=-0.024668606               pvth0=3.2106572e-014             pk2=4.8414672e-014 pminv=-2.3901559e-014            pvoff=-1.2740703e-013            peta0=7.1709773e-014 pu0=7.3539338e-015             pua=9.1733062e-023             pub=4.5866531e-031 puc=1.8515911e-022             pa0=-2.3697708e-012            pags=2.5481406e-014 pketa=-1.2995517e-013            wpclm=5.65625e-008               ppclm=-5.0962812e-013 ppdiblc2=1.0702191e-014             pkt1=-5.4065258e-028            pkt2=9.5689051e-014 pute=1.793891e-013              pua1=-1.4052486e-021            pub1=4.6138673e-030 puc1=-3.4141884e-022            pat=1.9539142e-008             wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.7 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.13199306 k2=0.0034018229               minv=-0.171365                  cit=0.0001 voff=-0.098606181               eta0=0.21595457                 etab=0.013821434 u0=0.044075903                ua=-1.3576389e-011            ub=3.0026215e-018 uc=3.5714311e-011             vsat=78486.111                  a0=6.9122396 ags=1.6671007                  keta=-0.015548611               pclm=1.8142361 pdiblc2=0.0066194444               tvoff=0.00130567                 ltvoff=3.51834e-009 wtvoff=1.03815e-009               ptvoff=-1.15415e-015              kt1=-0.18646875 kt2=-0.032801376               ute=-2.0482278                 ua1=5.4561632e-010 ub1=-4.1522642e-018            uc1=2.7273593e-012             at=153084.33 lvth0=-1.3700694e-009            lk2=6.4222005e-009             lvoff=-2.6031319e-010 leta0=-1.3456548e-007            lu0=-1.263204e-009             lua=-3.4251736e-017 lub=-3.9389496e-025            luc=-2.7711299e-018            la0=-1.7982161e-006 lags=-2.9113976e-007            lketa=-3.9732014e-008            lpclm=-3.4251736e-007 lpdiblc2=-3.8361944e-009            lkt1=1.8495937e-008             lkt2=3.321271e-008 lute=3.0141528e-007             lua1=6.3156091e-016             lub1=2.8641302e-025 luc1=-9.4324945e-017            lat=-0.13311252                letab=-6.9167956e-009 lvsat=0.0027401389               lcit=0                          wvth0=1.16625e-008 wk2=2.4133594e-008             wminv=-4.19985e-007              wvoff=-1.2544375e-008 weta0=-1.8334112e-007            wu0=-3.043875e-009             wua=7.84375e-017 wub=-5.7046875e-025            wuc=6.6097401e-017             wa0=-7.7126563e-006 wags=4.2421875e-007             wketa=-2.93125e-008              wpdiblc2=5.8625e-009 wkt1=3.509375e-008              wkt2=6.8352633e-008             wute=1.26925e-007 wua1=-3.5843437e-016            wub1=1.0768981e-024             wuc1=-2.4997118e-016 wat=-0.035928969               pvth0=7.398375e-015              pk2=-2.8206305e-014 pvoff=2.3428188e-015             peta0=1.7531683e-013             pu0=6.5845538e-015 pua=6.1653125e-023             pub=4.6239844e-031             puc=-6.9995779e-023 pa0=6.8126703e-012             pags=-4.6239844e-013            pketa=1.2330625e-014 wpclm=-5.65625e-007              ppclm=6.1653125e-013             ppdiblc2=-2.466125e-015 pkt1=-4.3157188e-014            pkt2=-1.0068726e-013            pute=-4.93225e-015 pua1=1.0394717e-022             pub1=-7.6079956e-032            puc1=3.5990548e-022 pat=3.9920398e-008             wetab=-6.8714281e-008            petab=1.2437285e-013 wvsat=0.002725                   pvsat=-4.93225e-009              wcit=0 pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.8 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.14288194 k2=0.016915964                minv=-0.44702111                cit=-0.0010545153 voff=-0.10410708                eta0=0.1609375                  etab=0.0023880556 u0=0.040239319                ua=-4.6776333e-011            ub=2.7755903e-018 uc=6.2007061e-011             vsat=81599.208                  a0=3.9190972 ags=1.9829861                  keta=-0.08636475                pclm=1.8548611 pdiblc2=0.0068006944               tvoff=-0.00114478                ltvoff=6.18933e-009 wtvoff=8.45551e-009               ptvoff=-9.23907e-015              kt1=-0.20338924 kt2=0.024415389                ute=-1.8393771                 ua1=1.5108502e-009 ub1=-5.6653264e-018            uc1=-2.6200832e-010            at=87361.08 lvth0=1.0498819e-008             lk2=-8.3082131e-009            lvoff=5.7356708e-009 leta0=-7.4596875e-008            lu0=2.9186718e-009             lua=1.9362033e-018 lub=-1.464309e-025             luc=-3.1430227e-017            la0=1.464309e-006 lags=-6.3545486e-007            lketa=3.7457578e-008             lpclm=-3.8679861e-007 lpdiblc2=-4.0337569e-009            lkt1=3.6939267e-008             lkt2=-2.9153564e-008 lute=7.3768021e-008             lua1=-4.2054403e-016            lub1=1.9356508e-024 luc1=1.9423695e-016             lat=-0.06147418                letab=5.5455869e-009 lvsat=-0.00065313708             lminv=3.0046516e-007             lcit=1.2584216e-009 wvth0=3.76125e-008               wk2=-3.9318675e-008            wminv=-6.052225e-007 wvoff=1.2821375e-007             weta0=-9.09375e-008              wu0=8.846125e-009 wua=1.50987e-016               wub=4.696875e-025              wuc=-1.394658e-016 wa0=8.803125e-006              wags=-6.84375e-007              wketa=3.578275e-008 wpdiblc2=6.79375e-009               wkt1=1.4045062e-007             wkt2=-7.273025e-008 wute=7.1141875e-007             wua1=5.5786062e-016             wub1=2.7983375e-024 wuc1=4.9172609e-016             wat=-0.037424894               pvth0=-2.0887125e-014 pk2=4.0956668e-014             pminv=2.0190888e-013             pvoff=-1.5108354e-013 peta0=7.4596875e-014             pu0=-6.3755462e-015            pua=-1.742583e-023 pub=-6.7137188e-031            puc=1.5406811e-022             pa0=-1.1189531e-011 pags=7.4596875e-013             pketa=-5.8623197e-014            wpclm=4.5625e-007 ppclm=-4.973125e-013             ppdiblc2=-3.4811875e-015            pkt1=-1.5799618e-013 pkt2=5.3093083e-014             pute=-6.4203044e-013            pua1=-8.9481438e-022 pub1=-1.9524489e-030            puc1=-4.4854454e-022            pat=4.1550957e-008 wetab=1.3715025e-007             petab=-1.0001949e-013            wvsat=-0.004637875 pvsat=3.0932837e-009             wcit=-2.0197275e-009            pcit=2.201503e-015 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.9 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.1233 k2=0.0075                     minv=-0.28585                   cit=0.0001 voff=-0.098363                  eta0=0.067493                   etab=0.01 u0=0.03995                    ua=3.5e-013                   ub=2.49e-018 uc=5.3288e-011                vsat=80000                      a0=4.525 ags=1.52                       keta=-0.00425                   pclm=1 pdiblc2=0.00185                    tvoff=0.004425                   ltvoff=0 wtvoff=-4.05e-010                 ptvoff=0                          kt1=-0.1725 kt2=-0.015521                  ute=-1.975                     ua1=5.327e-010 ub1=-2.709e-018                uc1=-5.478e-012                at=62500 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=-1.296e-008                wk2=2.7e-009 wminv=-2.0547e-007               wvoff=6.534e-010                 weta0=0 wu0=1.89e-009                  wua=2.97e-018                  wub=1.08e-025 wuc=-2.15028e-017              wa0=1.593e-006                 wags=-5.4e-007 wketa=-1.485e-008                wpdiblc2=2.7e-010                   wkt1=1.35e-008 wute=2.43e-007                  wua1=7.36668e-016               wub1=-6.3828e-025 wuc1=-3.82536e-017              wat=0.0135                     pvth0=0 pk2=0                          pvoff=0                          peta0=0 pu0=0                          pags=0                          ppdiblc2=0 wvsat=0                          pvsat=0                          wcit=0 pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.10 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.12478319 k2=0.006934375                minv=-0.28290246                cit=0.0001 voff=-0.098865778               eta0=0.081639407                etab=0.058360938 u0=0.038595768                ua=-7.1036806e-012            ub=2.4145833e-018 uc=5.4861192e-011             vsat=80000                      a0=4.5988832 ags=1.4659514                  keta=0.00366875                 pclm=0.98743056 pdiblc2=-0.00050048611             tvoff=0.00514498                 ltvoff=-6.487e-009 wtvoff=-1.37154e-009              ptvoff=8.70853e-015               kt1=-0.17312847 kt2=-0.020635664               ute=-1.9741704                 ua1=6.0054986e-010 ub1=-2.5752485e-018            uc1=2.6196573e-011             at=60098.105 lvth0=1.3363582e-008             lk2=5.0962812e-009             lvoff=4.5300278e-009 leta0=-1.2745913e-007            lu0=1.220163e-008              lua=6.7157662e-017 lub=6.7950417e-025             luc=-1.4174457e-017            la0=-6.6568758e-007 lags=4.8697799e-007             lketa=-7.1347937e-008            lpclm=1.1325069e-007 lpdiblc2=2.117788e-008              lkt1=5.6625347e-009             lkt2=4.6083123e-008 lute=-7.4745458e-009            lua1=-6.1132725e-016            lub1=-1.2051006e-024 luc1=-2.853879e-016             lat=0.021641075                letab=-4.3573205e-007 lvsat=0                          lminv=-2.6557288e-008            lcit=0 wvth0=-1.32315e-008              wk2=2.496375e-009              wminv=-2.0865334e-007 wvoff=4.7259e-009                weta0=-3.726066e-008             wu0=3.1022475e-009 wua=3.716625e-018              wub=2.166e-025                 wuc=-2.7989749e-017 wa0=2.2224727e-006             wags=-6.146625e-007             wketa=-1.2135e-008 wpdiblc2=2.238375e-009              wkt1=1.689375e-008              wkt2=5.5238372e-009 wute=2.291535e-007              wua1=7.1166285e-016             wub1=-7.1816887e-025 wuc1=-7.2162945e-017            wat=0.016993526                pvth0=2.446215e-015 pk2=1.8346612e-015             pminv=2.8681871e-014             pvoff=-3.6693225e-014 peta0=3.3571855e-013             pu0=-1.092235e-014             pua=-6.7270913e-024 pub=-9.78486e-031              puc=5.8447415e-023             pa0=-5.6715495e-012 pags=6.7270913e-013             pketa=-2.446215e-014             wpclm=-2.03625e-007 ppclm=1.8346612e-012             ppdiblc2=-1.7735059e-014            pkt1=-3.0577687e-014 pkt2=-4.9769773e-014            pute=1.2475697e-013             pua1=2.252964e-022 pub1=7.1979876e-031             puc1=3.055232e-022              pat=-3.1476671e-008 wetab=-8.7049687e-008            petab=7.8431768e-013             wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.11 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.10778681 k2=0.0077630208               minv=-0.297575                  cit=0.0011922708 voff=-0.079389278               eta0=-0.024780278               etab=-0.49136729 u0=0.043963903                ua=3e-011                     ub=2.7748611e-018 uc=4.7788307e-011             vsat=80000                      a0=2.4236681 ags=2.1967361                  keta=0.00171875                 pclm=-0.76666667 pdiblc2=0.018618056                tvoff=-0.00283102                ltvoff=7.94955e-009 wtvoff=8.48418e-009               ptvoff=-9.13033e-015              kt1=-0.18968056 kt2=0.036212273                ute=-2.4344347                 ua1=-1.1502866e-009 ub1=-2.5159729e-018            uc1=-2.4003129e-010            at=136366.77 lvth0=-1.7399882e-008            lk2=3.5964323e-009             lvoff=-3.0722437e-008 leta0=6.5160503e-008             lu0=2.485306e-009              lub=2.7401389e-026 luc=-1.3725356e-018            la0=3.2714518e-006             lags=-8.3574236e-007 lketa=-6.7818438e-008            lpclm=3.2881667e-006             lpdiblc2=-1.3426681e-008 lkt1=3.5621806e-008             lkt2=-5.6811642e-008            lute=8.2560385e-007 lua1=2.5576867e-015             lub1=-1.3123895e-024            luc1=1.9648454e-016 lat=-0.11640521                letab=5.5927605e-007             lvsat=0 lcit=-1.9770102e-009            wvth0=-3.190875e-008             wk2=1.6283437e-008 wminv=-1.92807e-007              wvoff=-4.71348e-008              weta0=2.499816e-007 wu0=-2.842275e-009             wub=-1.605e-025                wuc=4.4364208e-017 wa0=3.667725e-007              wags=-5.29125e-007              wketa=-6.039375e-008 wpdiblc2=-1.5735e-008               wkt1=4.0875e-008                wkt2=-5.5871934e-008 wute=8.220975e-007              wua1=2.6941909e-015             wub1=-1.8684263e-024 wuc1=1.869944e-016              wat=-0.0058373625              pvth0=3.6252037e-014 pk2=-2.3119922e-014            pvoff=5.7174642e-014             peta0=-1.8418994e-013 pu0=-1.6276425e-016            pub=-2.95935e-031              puc=-7.2513249e-023 pa0=-2.312732e-012             pags=5.1788625e-013             pketa=6.2886187e-014 wpclm=4.08e-006                  ppclm=-5.9187e-012               ppdiblc2=1.479675e-014 pkt1=-7.398375e-014             pkt2=6.1356573e-014             pute=-9.4847168e-013 pua1=-3.3630793e-021            pub1=2.8017646e-030             puc1=-1.6355159e-022 pat=9.8472371e-009             wetab=8.4062543e-007             petab=-8.9477427e-013 wvsat=0                          pvsat=0                          wcit=-1.9660875e-009 pcit=3.5586184e-015 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.12 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.13246944 k2=0.011388972                minv=-0.40418542                cit=-0.0043611278 voff=-0.072240972               eta0=-0.0045416667              etab=0.067924806 u0=0.050033917                ua=4.7763333e-011             ub=3.5806944e-018 uc=-1.6496971e-011            vsat=79022.611                  a0=11.457639 ags=1.1765278                  keta=-0.11733861                pclm=3.7708333 pdiblc2=0.00995                    tvoff=0.00489234                 ltvoff=-4.6891e-010 wtvoff=-2.41132e-009              ptvoff=2.74576e-015               kt1=-0.087548611 kt2=-0.11938245                ute=-1.0819486                 ua1=2.9816632e-009 ub1=-4.7592361e-018            uc1=2.6294189e-010             at=62357.097 lvth0=9.5041944e-009             lk2=-3.5585472e-010            lvoff=-3.851409e-008 leta0=4.3100417e-008             lu0=-4.1310092e-009            lua=-1.9362033e-017 lub=-8.5095694e-025            luc=6.8698417e-017             la0=-6.5755764e-006 lags=2.7628472e-007             lketa=6.1954086e-008             lpclm=-1.6577083e-006 lpdiblc2=-3.9785e-009               lkt1=-7.5702014e-008            lkt2=1.1278661e-007 lute=-6.4860601e-007            lua1=-1.9461385e-015            lub1=1.1327674e-024 luc1=-3.5175624e-016            lat=-0.035734666               letab=-5.0352338e-008 lvsat=0.0010653539               lminv=1.1620535e-007             lcit=4.0761943e-009 wvth0=1.887e-008                 wk2=-2.937009e-008             wminv=-6.8232675e-007 wvoff=7.085475e-008              weta0=2.06925e-007               wu0=-8.78415e-009 wua=-1.91844e-017              wub=-9.795e-025                wuc=1.8414585e-018 wa0=-4.76625e-006              wags=7.6725e-007                wketa=9.15357e-008 wpdiblc2=1.125e-009                 wkt1=-6.80625e-008              wkt2=1.8610586e-007 wute=-6.519525e-007             wua1=-2.0896027e-015            wub1=1.167375e-024 wuc1=-4.5318429e-016            wat=0.007582275                pvth0=-1.90968e-014 pk2=2.6642423e-014             pminv=5.3357653e-013             pvoff=-7.1433968e-014 peta0=-1.3725825e-013            pu0=6.3138795e-015             pua=2.0910996e-023 pub=5.96775e-031               puc=-2.6163452e-023            pa0=3.2822625e-012 pags=-8.951625e-013             pketa=-1.0271691e-013            wpclm=-2.9925e-006 ppclm=1.790325e-012              ppdiblc2=-3.58065e-015              pkt1=4.4758125e-014 pkt2=-2.0239923e-013            pute=6.5824283e-013             pua1=1.8512557e-021 pub1=-5.0725875e-031            puc1=5.3424318e-022             pat=-4.7801678e-009 wetab=1.91841e-008               petab=5.96775e-016               wvsat=0 pvsat=0                          wcit=3.932175e-009              pcit=-2.8704878e-015 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.13 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.14033571 k2=0.012766429                minv=-0.4761                    cit=0.0001 voff=-0.096329429               eta0=0.067493                   etab=0.013051357 u0=0.041477857                ua=-1.5145e-011               ub=2.7757143e-018 uc=2.1125857e-011             vsat=80000                      a0=7.2857143 ags=1.0574286                  keta=-0.024964286               pclm=1 pdiblc2=0.0021714286               tvoff=0.00405286                 ltvoff=0 wtvoff=-3.08571e-012              ptvoff=0                          kt1=-0.13682143 kt2=-0.015521                  ute=-1.7142857                 ua1=1.5591571e-009 ub1=-3.8617143e-018            uc1=-3.8385143e-011            at=75000 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=5.4385714e-009             wk2=-2.9877429e-009 wvoff=-1.5428571e-009            weta0=0                          wu0=2.3991429e-010 wua=1.97046e-017               wub=-2.0057143e-025            wuc=1.3232314e-017 wa0=-1.3885714e-006            wags=-4.0422857e-008            wketa=7.5214286e-009 wpdiblc2=-7.7142857e-011            wkt1=-2.5032857e-008            wute=-3.8571429e-008 wua1=-3.7190571e-016            wub1=6.0665143e-025             wuc1=-2.7138857e-018 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wetab=-3.2954657e-009            wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.14 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.14344396 k2=0.013628333                minv=-0.4761                    cit=0.0001 voff=-0.097953042               eta0=0.042028419                etab=-0.028573274 u0=0.041150369                ua=-2.4698317e-011            ub=2.811627e-018 uc=1.8244874e-011             vsat=80000                      a0=8.034451 ags=0.93288333                 keta=-0.018167808               pclm=0.76297619 pdiblc2=0.0022540278               tvoff=0.00381828                 ltvoff=2.11358e-009 wtvoff=6.12986e-011               ptvoff=-5.80102e-016              kt1=-0.13386761 kt2=-0.021283821               ute=-1.7207464                 ua1=1.6314709e-009 ub1=-3.8484589e-018            uc1=-3.3831269e-011            at=75529.928 lvth0=2.8005279e-008             lk2=-7.7657619e-009            lvoff=1.4628754e-008 leta0=2.2943588e-007             lu0=2.950666e-009              lua=8.6075381e-017 lub=-3.2357341e-025            luc=2.5957658e-017             la0=-6.7461174e-006 lags=1.1221526e-006             lketa=-6.1236268e-008            lpclm=2.1355845e-006 lpdiblc2=-7.4421885e-010            lkt1=-2.6613913e-008            lkt2=5.1923017e-008 lute=5.8210857e-008             lua1=-6.5154742e-016            lub1=-1.1943095e-025 luc1=-4.1030403e-017            lat=-0.0047746493              letab=3.7503793e-007 lvsat=0                          lcit=0                          wvth0=6.922125e-009 wk2=-4.7331e-009               wvoff=3.740145e-009              weta0=5.5192071e-009 wu0=3.4327821e-010             wua=2.2718832e-017             wub=-2.1220714e-025 wuc=1.1555874e-017             wa0=-1.4879404e-006            wags=-3.8949e-008 wketa=1.1448482e-008             wpdiblc2=-7.365e-010                wkt1=-2.5507982e-008 wkt2=6.2238466e-009             wute=-4.4544429e-008            wua1=-4.0173193e-016 wub1=6.5689832e-025             wuc1=-7.3328764e-018            wat=0.0003271575 pvth0=-1.3366818e-014            pk2=1.5725668e-014             pvoff=-4.7599849e-014 peta0=-4.9728056e-014            pu0=-9.31309e-016              pua=-2.7158228e-023 pub=1.0483779e-031             puc=1.5104731e-023             pa0=8.9531469e-013 pags=-1.3279453e-014            pketa=-3.5382753e-014            wpclm=3.8785714e-008 ppclm=-3.4945929e-013            ppdiblc2=5.9408079e-015             pkt1=4.2808763e-015 pkt2=-5.6076858e-014            pute=5.381673e-014              pua1=2.6873419e-022 pub1=-4.527245e-031             puc1=4.1617106e-023             pat=-2.9476891e-009 wetab=6.8392608e-009             petab=-9.1313886e-014            wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.15 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.14760873 k2=0.027789459                minv=-0.4761                    cit=-0.00082390476 voff=-0.12172654                eta0=0.27400817                 etab=0.40296346 u0=0.041542643                ua=4.3790476e-012             ub=2.8216607e-018 uc=9.2651253e-011             vsat=81297.619                  a0=3.6695778 ags=1.4468849                  keta=-0.064543651               pclm=3.9109127 pdiblc2=-0.004282121               tvoff=0.00521724                 ltvoff=-4.18537e-010 wtvoff=-2.07931e-010              ptvoff=-9.27968e-017              kt1=-0.14986905 kt2=0.007634878                ute=-1.7175875                 ua1=1.5074547e-009 ub1=-4.532023e-018             uc1=-8.1053115e-011            at=135534.13 lvth0=3.5543516e-008             lk2=-3.33974e-008              lvoff=5.7658785e-008 leta0=-1.9044748e-007            lu0=2.2406507e-009             lua=3.3445352e-017 lub=-3.4173446e-025            luc=-1.0871789e-016            la0=1.1543031e-006 lags=1.9180972e-007             lketa=2.2704008e-008             lpclm=-3.5621806e-006 lpdiblc2=1.1086211e-008             lkt1=2.3486905e-009             lkt2=-4.1982842e-010 lute=5.2493232e-008             lua1=-4.2707805e-016            lub1=1.1178201e-024 luc1=4.4441138e-017             lat=-0.11338225                letab=-4.0604357e-007 lvsat=-0.0023486905              lcit=1.6722676e-009             wvth0=1.1098929e-008 wk2=-5.3451161e-009            wvoff=-1.4105571e-009            weta0=-7.2709929e-008 wu0=-2.2731429e-010            wua=2.7670629e-017             wub=-2.1104357e-025 wuc=-4.0877729e-018            wa0=-9.7881e-007               wags=2.8071429e-007 wketa=1.1169643e-008             wpdiblc2=8.9971907e-009             wkt1=-2.1214286e-009 wkt2=-2.5008348e-008            wute=4.79025e-008               wua1=-1.7616975e-016 wub1=3.0890786e-025             wuc1=1.5297964e-017             wat=-0.0049381071 pvth0=-2.0926832e-014            pk2=1.6833417e-014             pvoff=-3.8277078e-014 peta0=9.1866679e-014             pu0=1.0146343e-016             pua=-3.6120981e-023 pub=1.0273172e-031             puc=4.3419731e-023             pa0=-2.6211386e-014 pags=-5.9187e-013               pketa=-3.4878054e-014            wpclm=-9.7178571e-007 ppclm=1.479675e-012              ppdiblc2=-1.1677172e-014            pkt1=-3.8048786e-014 pkt2=4.534147e-016              pute=-1.1351221e-013            pua1=-1.3953335e-022 pub1=1.7713824e-031             puc1=6.5528464e-025             pat=6.5824399e-009 wetab=-1.2525179e-007            petab=1.4777092e-013             wvsat=-0.0014014286 pvsat=2.5365857e-009             wcit=2.1138214e-010             pcit=-3.8260168e-016 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na18_mac.16 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.095765079 k2=-0.03964004                minv=-1.1083901                 cit=-0.00065133809 voff=0.081284921                eta0=0.16330556                 etab=0.059083575 u0=0.043725167                ua=5.9813333e-011             ub=3.051877e-018 uc=-6.376962e-011             vsat=76018.921                  a0=10.247024 ags=2.3325794                  keta=0.017119048                pclm=-0.081349206 pdiblc2=0.016091623                tvoff=0.00485724                 ltvoff=-2.61444e-011 wtvoff=-2.37341e-009              ptvoff=2.26757e-015               kt1=-0.11411111 kt2=0.076537722                ute=-1.5808147                 ua1=1.8498085e-009 ub1=-4.9514365e-018            uc1=-1.5588913e-010            at=74673.516 lvth0=-2.0966063e-008            lk2=4.0100754e-008             lvoff=-1.6362371e-007 leta0=-6.9781627e-008            lu0=-1.3830024e-010            lua=-2.6978019e-017 lub=-5.926702e-025             luc=6.1780863e-017             la0=-6.0151131e-006 lags=-7.7359722e-007            lketa=-6.6308333e-008            lpclm=7.8938492e-007 lpdiblc2=-1.1121171e-008            lkt1=-3.662746e-008             lkt2=-7.5523929e-008 lute=-9.6589139e-008            lua1=-8.002437e-016             lub1=1.5749808e-024 luc1=1.2601239e-016             lat=-0.047044184               letab=-3.121449e-008 lvsat=0.0034050908               lminv=6.8919619e-007             lcit=1.4841699e-009 wvth0=-2.0770714e-008            wk2=2.5741243e-008             wminv=7.8214286e-008 wvoff=-9.4953214e-008            weta0=2.565e-008                 wu0=-1.9707e-009 wua=-3.21984e-017              wub=-4.0837714e-025            wuc=5.2895919e-017 wa0=-3.4587857e-006            wags=-4.8128571e-007            wketa=-5.3678571e-008 wpdiblc2=-5.5079529e-009            wkt1=-3.9375e-008               wkt2=-2.5487925e-008 wute=-1.1317714e-007            wua1=-8.6719971e-016            wub1=1.3749514e-024 wuc1=-8.46786e-019              wat=-0.0057194571              pvth0=1.3811079e-014 pk2=-1.7050714e-014            pminv=-8.5253571e-014            pvoff=6.3684418e-014 peta0=-1.5345643e-014            pu0=2.0017539e-015             pua=2.9136261e-023 pub=3.1782531e-031             puc=-1.8692494e-023            pa0=2.6769621e-012 pags=2.3871e-013                pketa=3.58065e-014               wpclm=1.1678571e-006 ppclm=-8.5253571e-013            ppdiblc2=4.1334342e-015             pkt1=2.5576071e-015 pkt2=9.7615339e-016             pute=6.20646e-014               pua1=6.1368931e-022 pub1=-9.8484926e-031            puc1=1.8253063e-023             pat=7.4341114e-009 wetab=2.8732629e-008             petab=-2.0072101e-014            wvsat=0.0032439857 pvsat=-2.5269159e-009            wcit=-7.4397857e-011            pcit=-7.1101479e-017 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.prot
.option tmiflag=2.01 modmonte=1 tmipath='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.option etmiUsrInput='/proj/db40/a0/staff/jcorn/rbdata/cad/models/spice/FOUNDRY/TMI/model_card/cln45gs_1d2_1d8_ud15_lk_v2d0_2_tmi_v1d0_dir'
.unprot
.model nch_na18ud15_mac.global nmos ( modelid=16                         level=54                         version=4.5 binunit=2                          paramchk=1                          mobmod=0 capmod=2                          igcmod=0                          igbmod=0 diomod=1                          rdsmod=0                          rbodymod=0 rgatemod='1*rgflag_na18ud15'        permod=1                          acnqsmod=0 trnqsmod=0                          tempmod=0                          tnom=25 toxe=3.36e-009                  toxm=3.36e-009                  dtox=1.9844e-010 epsrox=3.9                        wint=0                          lint=0 ll=0                          wl=0                          lln=1 wln=1                          lw=0                          ww=0 lwn=1                          wwn=1                          lwl=0 wwl=0                          llc=0                          wlc=0 lwc=0                          wwc=0                          lwlc=0 wwlc=0                          xl=1e-008                     xw=0 dlc=3.542614e-008              dwc=0                          xpart=1 toxref=3e-009                     dlcig=2.5e-009                   k1=0.054 k3=-8.2825                    k3b=-4.2795                    w0=0 dvt0=0.0050825                  dvt1=45.501                     dvt2=0.185 dvt0w=0                          dvt1w=0                          dvt2w=0 dsub=0.062479                   voffl=-5e-009                    dvtp0=0 dvtp1=4                          lpe0=-4.24e-007                 lpeb=-1e-007 xj=6.7e-008                   ngate=3e+021                     ndep=1e+017 nsd=1e+020                     phin=0.19                       cdsc=0 cdscb=0                          cdscd=0                          nfactor=0.53 ud=0                          lud=0                          wud=0 pud=0                          a1=0                          a2=1 b0=0                          b1=0                          dwg=0 dwb=0                          pdiblc1=0                          pdiblcb=0 drout=0.56                       pvag=0.3                        delta=0.01 pscbe1=9.264e+008                 pscbe2=1e-020                     fprout=100 pdits=0                          pditsd=0                          pditsl=0 rsh=18.0                       rdsw=217.15                     prwg=0 prwb=0                          wr=1                          alpha0=0 alpha1=0.00035                    beta0=7                          agidl=1.4314e-011 bgidl=2.3e+009                   cgidl=0.5                        egidl=0.8 aigbacc=0.01238                    bigbacc=0.006109                   cigbacc=0.2809 nigbacc=4.05                       aigbinv=0.0111                     bigbinv=0.000949 cigbinv=0.006                      eigbinv=1.1                        nigbinv=1 aigc=0.009898                   bigc=0.001383                   cigc=1.515e-005 aigsd=0.0086                     bigsd=0.0004353                  cigsd=3.925e-020 nigc=1                          poxedge=1                          pigcd=1.672 ntox=1                          xrcrg1=12                         xrcrg2=1 vfbsdoff=0                          lvfbsdoff=0                          wvfbsdoff=0 pvfbsdoff=0                          cgso=4.925043e-011              cgdo=4.925043e-011 cgbo=0                          cgdl=3.247859e-010              cgsl=3.247859e-010 clc=0                          cle=0.6                        cf='8.050e-11+7.81e-11*ccoflag_na18ud15' ckappas=0.6                        ckappad=0.6                        acde=0.3 moin=16.193                     noff=3.9                        voffcv=-0.004675 kt1l=0                          prt=0                          fnoimod=1.000000e+00 tnoimod=0                          em=1.300000e+06               ef=1.050000e+00 noia=0                          noib=0                          noic=0 lintnoi=-1.000000e-07              jss=1.60e-06                   jsd=1.60e-06 jsws=1.57e-12                   jswd=1.57e-12                   jswgs=1.57e-12 jswgd=1.57e-12                   njs=1.02                       njd=1.02 ijthsfwd=0.01                       ijthdfwd=0.01                       ijthsrev=0.01 ijthdrev=0.01                       bvs=19.65                      bvd=19.65 xjbvs=1                          xjbvd=1                          jtsswgs=1.6e-010 jtsswgd=1.6e-010                   njtsswg=20                         xtsswgs=0.69066 xtsswgd=0.69066                    tnjtsswg=1                          vtsswgs=10 vtsswgd=10                         pbs=0.512                      pbd=0.512 cjs=0.000161                   cjd=0.000161                   mjs=0.292 mjd=0.292                      pbsws=0.3                        pbswd=0.3 cjsws=2.08e-010                  cjswd=2.08e-010                  mjsws=0.039 mjswd=0.039                      pbswgs=0.791                      pbswgd=0.791 cjswgs=1.62e-010                  cjswgd=1.62e-010                  mjswgs=0.385 mjswgd=0.385                      tpb=0.0014                     tcj=0.0012 tpbsw=0.0013                     tcjsw=0.00034                    tpbswg=0.0022 tcjswg=0.0015                     xtis=3                          xtid=3 dmcg=6.7e-008                   dmci=6.7e-008                   dmdg=0 dmcgt=0                          dwj=0                          xgw=0 xgl=2.64e-09                   rshg=16.42                      gbmin=1e-012 rbpb=50                         rbpd=50                         rbps=50 rbdb=50                         rbsb=50                         ngcon=1 lnfactor=0                          pnfactor=0                          rdw=0 rsw=0                          wnfactor=0 tmimodel=1 tmi_ver=101011.200002 tmi_ver_inst=0.1                       tmi_ver_weflef=0.1                     tmi_ver_nrsd=0.2 tmi_ver_adaspdps=0.1                   tmi_ver_rdr=0.0                        tmi_ver_mclib=0.1 tmi_ver_mcratio=0.1                    tmi_ver_mcglobal=0.2                   tmi_ver_mclocal=0.2 tmi_ver_mcdelta=0.3                    tmi_ver_mccorsum=0.2                   tmi_ver_iboff=0.0 tmi_ver_lod=0.2                        tmi_ver_pse=0.2                        tmi_ver_cesl=0.1 tmi_ver_ose=0.2                        tmi_ver_wpe=0.1                        tmi_ver_cf=0.1 tmi_ver_tnoi=0.7 sigma_factor='sigma_factor_na18ud15' ccoflag='ccoflag_na18ud15' rcoflag='rcoflag_na18ud15' rgflag='rgflag_na18ud15' mismatchflag='mismatchflag_mos_na18ud15' globalflag='globalflag_mos_na18ud15' totalflag='totalflag_mos_na18ud15' global_factor='global_factor_na18ud15' local_factor='local_factor_na18ud15' sigma_factor_flicker='sigma_factor_flicker_na18ud15' noiseflag='noiseflagn_na18ud15' noiseflag_mc='noiseflagn_na18ud15_mc' delvto=0 mulu0=1 dlc_fmt=2 par1_io='par1_io' par2_io='par2_io' par3_io='par3_io' par4_io='par4_io' par5_io='par5_io' par6_io='par6_io' par7_io='par7_io' par8_io='par8_io' par9_io='par9_io' par10_io='par10_io' par11_io='par11_io' par12_io='par12_io' par13_io='par13_io' par14_io='par14_io' par15_io='par15_io' par16_io='par16_io' par17_io='par17_io' par18_io='par18_io' par19_io='par19_io' par20_io='par20_io' w1_io='2.0857*0.40825' w2_io='0.67082*-0.40825' w3_io='0.54772*0.26807' w4_io='0.54772*-0.6902' w5_io='0.54772*-0.32981' w6_io='0.54772*0.098267' tox_c='toxn_na18ud15'            dxl_c='dxln_na18ud15'            dxw_c='dxwn_na18ud15' cj_c='cjn_na18ud15'             cjsw_c='cjswn_na18ud15'           cjswg_c='cjswgn_na18ud15' cgo_c='cgon_na18ud15'            cgl_c='cgln_na18ud15'            ddlc_c='ddlcn_na18ud15' dvth_c='dvthn_na18ud15'           dlvth_c='dlvthn_na18ud15'          dwvth_c='dwvthn_na18ud15' dpvth_c='dpvthn_na18ud15'          cf_c='cfn_na18ud15'             du0_c='du0n_na18ud15' dlu0_c='dlu0n_na18ud15'           dwu0_c='dwu0n_na18ud15'           dpu0_c='dpu0n_na18ud15' dvsat_c='dvsatn_na18ud15'          dlvsat_c='dlvsatn_na18ud15'         dwvsat_c='dwvsatn_na18ud15' dpvsat_c='dpvsatn_na18ud15'         dk2_c='dk2n_na18ud15'            drdsw_c='drdswn_na18ud15' dvoff_c='dvoffn_na18ud15'          dlvoff_c='dlvoffn_na18ud15'         dwvoff_c='dwvoffn_na18ud15' dpvoff_c='dpvoffn_na18ud15'         dpdiblc2_c='dpdiblc2n_na18ud15'       dlpdiblc2_c='dlpdiblc2n_na18ud15' dwpdiblc2_c='dwpdiblc2n_na18ud15'      dppdiblc2_c='dppdiblc2n_na18ud15'      dags_c='dagsn_na18ud15' dlags_c='dlagsn_na18ud15'          dwags_c='dwagsn_na18ud15'          dpags_c='dpagsn_na18ud15' dnfactor_c='dnfactorn_na18ud15'       dlnfactor_c='dlnfactorn_na18ud15'      dwnfactor_c='dwnfactorn_na18ud15' dpnfactor_c='dpnfactorn_na18ud15'      dcit_c='dcitn_na18ud15'           dlcit_c='dlcitn_na18ud15' dwcit_c='dwcitn_na18ud15'          dpcit_c='dpcitn_na18ud15'          deta0_c='deta0n_na18ud15' dleta0_c='dleta0n_na18ud15'         dweta0_c='dweta0n_na18ud15'         dpeta0_c='dpeta0n_na18ud15' dub1_c='dub1n_na18ud15'           dlk2_c='dlk2n_na18ud15'           dwk2_c='dwk2n_na18ud15' dpk2_c='dpk2n_na18ud15'           dkt1_c='dkt1n_na18ud15'           dlkt2_c='dlkt2n_na18ud15' dla0_c='dla0n_na18ud15'           dwa0_c='dwa0n_na18ud15'           dluc_c='dlucn_na18ud15' dlketa_c='dlketan_na18ud15'         monte_flag_c='monte_flagn_na18ud15'    c1f_c='c1fn_na18ud15' c2f_c='c2fn_na18ud15'            c3f_c='c3fn_na18ud15' global_mc='global_mc_flag_na18ud15' tox_g='toxn_na18ud15_ms_global'  dxl_g='dxln_na18ud15_ms_global' dxw_g='dxwn_na18ud15_ms_global'  cj_g='cjn_na18ud15_ms_global' cjsw_g='cjswn_na18ud15_ms_global' cjswg_g='cjswgn_na18ud15_ms_global' cgo_g='cgon_na18ud15_ms_global'  cgl_g='cgln_na18ud15_ms_global' dvth_g='dvthn_na18ud15_ms_global' dlvth_g='dlvthn_na18ud15_ms_global' dwvth_g='dwvthn_na18ud15_ms_global'                                        dpvth_g='dpvthn_na18ud15_ms_global' cf_g='cfn_na18ud15_ms_global'   du0_g='du0n_na18ud15_ms_global' dlu0_g='dlu0n_na18ud15_ms_global' dwu0_g='dwu0n_na18ud15_ms_global' dpu0_g='dpu0n_na18ud15_ms_global' dvsat_g='dvsatn_na18ud15_ms_global' dlvsat_g='dlvsatn_na18ud15_ms_global'                                       dwvsat_g='dwvsatn_na18ud15_ms_global' dpvsat_g='dpvsatn_na18ud15_ms_global'                                       dk2_g='dk2n_na18ud15_ms_global' dlvoff_g='dlvoffn_na18ud15_ms_global'                                       dppdiblc2_g='dppdiblc2n_na18ud15_ms_global' dags_g='dagsn_na18ud15_ms_global' dwags_g='dwagsn_na18ud15_ms_global' deta0_g='deta0n_na18ud15_ms_global'                                        dlk2_g='dlk2n_na18ud15_ms_global' dwk2_g='dwk2n_na18ud15_ms_global' dpk2_g='dpk2n_na18ud15_ms_global' dkt1_g='dkt1n_na18ud15_ms_global' dlkt2_g='dlkt2n_na18ud15_ms_global' dla0_g='dla0n_na18ud15_ms_global' dwa0_g='dwa0n_na18ud15_ms_global' dluc_g='dlucn_na18ud15_ms_global' dlketa_g='dlketan_na18ud15_ms_global' monte_flag_g='monte_flagn_na18ud15_ms_global'                                  ddlc_g='ddlcn_na18ud15_ms_global' weight1=-3.1983125 weight2=1.5975625 weight3=-1.038375 weight4=-0.625 weight5=-0.4297125 tox_1=1.2526e-011 tox_2=-2.6961e-011 tox_3=-1.0998e-012 tox_4=9.4257e-011 tox_5=4.0716e-012 dxl_1=7.5174e-010 dxl_2=-1.618e-009 dxl_3=-6.6005e-011 dxl_4=-5.6569e-009 dxl_5=2.4436e-010 dxw_1=-1.2161e-009 dxw_2=-2.3698e-009 dxw_3=-1.3015e-009 dxw_4=-2.1115e-024 dxw_5=-1.1627e-008 cj_1=1.0896e-006 cj_2=-1.1204e-007 cj_3=4.5396e-007 cj_4=2.0024e-021 cj_5=-1.431e-007 cjsw_1=1.4077e-012 cjsw_2=-1.4475e-013 cjsw_3=5.8648e-013 cjsw_4=-2.9972e-028 cjsw_5=-1.8487e-013 cjswg_1=1.0964e-012 cjswg_2=-1.1274e-013 cjswg_3=4.5678e-013 cjswg_4=5.2561e-028 cjswg_5=-1.4399e-013 cgo_1=-3.3333e-013 cgo_2=3.4274e-014 cgo_3=-1.3887e-013 cgo_4=4.3203e-028 cgo_5=4.3775e-014 cgl_1=-2.1982e-012 cgl_2=2.2602e-013 cgl_3=-9.1577e-013 cgl_4=3.2719e-027 cgl_5=2.8868e-013 dvth_1=0.006065 dvth_2=0.0034522 dvth_3=0.0032314 dvth_4=-3.8046e-018 dvth_5=-0.0016707 dlvth_1=1.3793e-009 dlvth_2=8.4963e-010 dlvth_3=5.4735e-010 dlvth_4=1.1923e-025 dlvth_5=-3.7158e-010 dwvth_1=3.7255e-010 dwvth_2=1.5998e-010 dwvth_3=1.4975e-010 dwvth_4=4.9101e-025 dwvth_5=-8.7014e-011 dpvth_1=4.8676e-017 dpvth_2=2.0468e-016 dpvth_3=-9.0892e-017 dpvth_4=-9.9193e-033 dpvth_5=-3.4886e-017 cf_1=-5.4482e-013 cf_2=5.6021e-014 cf_3=-2.2698e-013 cf_4=1.0968e-027 cf_5=7.155e-014 du0_1=4.8192e-005 du0_2=0.00047724 du0_3=0.00013197 du0_4=-1.5639e-019 du0_5=-0.00011294 dlu0_1=-1.7706e-011 dlu0_2=1.1738e-010 dlu0_3=2.1062e-011 dlu0_4=5.9835e-027 dlu0_5=-2.3406e-011 dwu0_1=3.0143e-013 dwu0_2=7.9941e-011 dwu0_3=1.5712e-013 dwu0_4=-1.9145e-026 dwu0_5=-1.8178e-011 dpu0_1=-1.2201e-017 dpu0_2=1.0069e-016 dpu0_3=-2.1616e-018 dpu0_4=3.3721e-032 dpu0_5=-2.0657e-017 dvsat_1=-966.86 dvsat_2=99.417 dvsat_3=-402.8 dvsat_4=-1.7393e-012 dvsat_5=126.97 dlvsat_1=0.00054684 dlvsat_2=-7.7595e-005 dlvsat_3=0.00042603 dlvsat_4=-5.1274e-019 dlvsat_5=-8.9805e-005 dwvsat_1=-0.00024778 dwvsat_2=1.1234e-005 dwvsat_3=2.8912e-005 dwvsat_4=-5.4722e-020 dwvsat_5=2.0547e-005 dpvsat_1=1.0777e-010 dpvsat_2=4.7294e-012 dpvsat_3=-1.0178e-010 dpvsat_4=1.3419e-025 dpvsat_5=-8.4078e-013 dk2_1=0.00013668 dk2_2=-1.7758e-005 dk2_3=9.13e-005 dk2_4=3.0668e-020 dk2_5=-2.1068e-005 dlvoff_1=-2.1765e-010 dlvoff_2=-3.4598e-011 dlvoff_3=4.3789e-010 dlvoff_4=2.7605e-025 dlvoff_5=-1.9391e-011 dppdiblc2_1=4.2274e-018 dppdiblc2_2=-1.8591e-018 dppdiblc2_3=1.4975e-017 dppdiblc2_4=-7.1959e-033 dppdiblc2_5=-1.7545e-018 dags_1=-0.002906 dags_2=0.00062643 dags_3=-0.0042499 dags_4=-3.596e-018 dags_5=0.00065749 dwags_1=1.39e-009 dwags_2=-5.7462e-011 dwags_3=-2.1375e-010 dwags_4=-1.0871e-024 dwags_5=-1.1059e-010 deta0_1=-0.0004502 deta0_2=4.4867e-005 deta0_3=-0.00017434 deta0_4=2.7218e-019 deta0_5=5.7923e-005 dlk2_1=4.5329e-011 dlk2_2=-3.8768e-013 dlk2_3=-2.0758e-011 dlk2_4=-5.0997e-026 dlk2_5=-2.3549e-012 dwk2_1=4.2316e-011 dwk2_2=4.1955e-012 dwk2_3=-6.1655e-011 dwk2_4=1.5331e-026 dwk2_5=1.6389e-012 dpk2_1=1.4503e-016 dpk2_2=-1.4913e-017 dpk2_3=6.042e-017 dpk2_4=1.3354e-031 dpk2_5=-1.9046e-017 dkt1_1=-0.0022058 dkt1_2=0.00015559 dkt1_3=-0.00025824 dkt1_4=1.1147e-018 dkt1_5=0.00022971 dlkt2_1=1.6324e-011 dlkt2_2=2.5948e-012 dlkt2_3=-3.2842e-011 dlkt2_4=7.5187e-027 dlkt2_5=1.4543e-012 dla0_1=7.8562e-008 dla0_2=-5.2293e-009 dla0_3=6.3016e-009 dla0_4=1.6764e-022 dla0_5=-7.9187e-009 dwa0_1=-1.783e-008 dwa0_2=-3.0324e-010 dwa0_3=1.2393e-008 dwa0_4=3.754e-023 dwa0_5=5.4259e-010 dluc_1=5.4412e-019 dluc_2=8.6494e-020 dluc_3=-1.0947e-018 dluc_4=7.0457e-034 dluc_5=4.8477e-020 dlketa_1=-2.7206e-010 dlketa_2=-4.3247e-011 dlketa_3=5.4736e-010 dlketa_4=2.4041e-026 dlketa_5=-2.4239e-011 monte_flag_1=0.0939675 monte_flag_2=-0.20225 monte_flag_3=-0.00825062 monte_flag_4=-0.707113 monte_flag_5=0.030545 sigma_local=1                          a_1=1 b_1=0                          c_1=0                          d_1=0 e_1_1=0                          e_1_2=0                          f_1_1=0 f_1_2=0                          g_1_1=0                          g_1_2=0 a_2=1                          b_2=0                          c_2=0 d_2=0                          a_3=1                          b_3=0 c_3=0                          d_3=0                          e_3_1=0 e_3_2=0                          f_3_1=0                          f_3_2=0 g_3_1=0                          g_3_2=0                          a_4=0.999982526 b_4=-4.20e-05                  c_4=-1.11e-04                  d_4=-1.04e-03 e_4_1=0                          e_4_2=0                          f_4_1=0 f_4_2=0                          g_4_1=5.0e-06                    g_4_2=1.04988e-08 a_5=1                          b_5=0                          c_5=0 d_5=0                          e_5_1=0                          e_5_2=0 f_5_1=0                          f_5_2=0                          g_5_1=0 g_5_2=0                          sigma_global=1 plo_tox='plo_tox'                  plo_dxl='plo_dxl' plo_dxw='plo_dxw'                  parl1='parl1'                    parl2='parl2' mis_a_1=0.00185                    mis_a_2=-0.015                     mis_a_3=-0.035 mis_b_1=0.0010                     mis_b_2=0.16                       mis_b_3=0.01 mis_c_1=1                          mis_c_2=0                          mis_c_3=0 mis_d_1=0.002                      mis_d_2=0                          mis_d_3=0 mis_e_1=0.0017                     mis_e_2=0                          mis_e_3=0.23 e_limit1=0.1                        e_limit2=2                          avtgm_min=0 d=0 xw0=0                          xl0=1e-8 co_enod=0.027                      co_size=0.054                      co_pitch=0.126 co_rc=52                         co_rsd=18.0                       bidirectionflag=1 designflag=1 cf0=8.050e-11                  cco=7.81e-11 noimod=1                          noic2='2.236'                    noic3='0.8' noiareac='0.81*9.5e-6*10e-6'        noic1=2.718 saref0=0.533e-6             sbref0=0.533e-6 samax=10e-6               sbmax=10e-6 samin=0.135e-6            sbmin=0.135e-6 rllodflag=0                   lreflod=1e-6                llodref=0.1 lod_clamp=-1e90 wlod0=1e-8 ku00=-3.0e-8             lku00=4e-6             wku00=0e-6 pku00=0.04e-11            tku00=0.8              llodku00=1 wlodku00=1                   kvsat0=0 kvth00=18.5e-9             lkvth00=14.0e-7          wkvth00=1.5e-6 pkvth00=0e-13               llodvth0=1                wlodvth0=1 stk20=7.5e-10             lodk20=1                steta00=-1.4e-9 lodeta00=1 wlod00=0 ku000=0e-8               lku000=0e-6               wku000=0e-6       		pku000=0.00e-11 llodku000=1                  wlodku000=1 kvth000=0e-8               lkvth000=-0e-15             wkvth000=-0e-15     		pkvth000=0 llodvth00=1                  wlodvth00=1                  steta000=-0e-9 stk200=0                  lodk200=1 lodeta000=1 wlod1=0                   llod1=0 ku01=0                   lku01=0                wku01=0 pku01=0                   llodku01=1 wlodku01=1                   kvsat1=0 kvth01=0                   lkvth01=0                wkvth01=0 pkvth01=0                   llodvth1=1                wlodvth1=1 steta01=0                   lodeta01=1 stk21=0                   lodk21=1 wlod2=0 ku02=0                   lku02=0                wku02=0 pku02=0                   tku02=0                llodku02=1 wlodku02=1                   kvsat2=1 kvth02=0                   lkvth02=0                wkvth02=0 pkvth02=0                   llodvth2=1                wlodvth2=1 stk22=0                   lodk22=1                steta02=0 lodeta02=1 wlod02=0 ku002=0                   lku002=0                   wku002=0                pku002=0 llodku002=1                   wlodku002=1 kvth002=0                   lkvth002=0                   wkvth002=0         		pkvth002=0 llodvth02=1                   wlodvth02=1                   steta002=0 stk202=0                   lodk202=1 lodeta002=1 wlod3=0 ku03=0                   lku03=0                wku03=0 pku03=0                   tku03=0                llodku03=1 wlodku03=1                   kvsat3=0 kvth03=0                   lkvth03=0                wkvth03=0 pkvth03=0                   llodvth3=1                wlodvth3=1 stk23=0                   lodk23=1                steta03=0 lodeta03=1 wlod03=0 ku003=0.0e-2              lku003=-0.0e-8              wku003=0         		pku003=0 llodku003=1                   wlodku003=1 kvth003=0                   lkvth003=0                   wkvth003=0         		pkvth003=0 llodvth03=1                   wlodvth03=1                   steta003=0 stk203=0                   lodk203=1 lodeta003=1 sa_b=5.33e-7             sa_b1=1.35e-7             dpdbinflag=0 w_b=9e-7                w_b1=5.4e-7 sparef=1.98e-7             spamax=1.6e-6              spamin=1.98e-7 kvth0dpc=0.00                wkvth0dpc=0.0e-8              wdpckvth0=1 lkvth0dpc=0.0e-8              ldpckvth0=1                   pkvth0dpc=0.0e-15 ku0dpc=0.00                wku0dpc=0.0e-8              wdpcku0=1 lku0dpc=0.0e-8              ldpcku0=1                   pku0dpc=0.0e-14 keta0dpc=0.000               wketa0dpc=0e-9                wdpcketa0=1 kvsatdpc=0.00                wdpc=0 kvth0dpc_b1=-0.000            kvth0dpc_b2=-0.000            dpcbinflg=0 ku0dpc_b1=0                 ku0dpc_b2=0 keta0dpc_b1=0                  keta0dpc_b2=0 kvth0dpl=0.05                wkvth0dpl=0.0e-8              wdplkvth0=1 lkvth0dpl=1.5e-6              ldplkvth0=0.8                 pkvth0dpl=0.0e-19 ku0dpl=0.20                wku0dpl=-3e-8               wdplku0=1 lku0dpl=6e-6                ldplku0=0.8                 pku0dpl=0.0e-11 keta0dpl=0                   wketa0dpl=0e-7                wdplketa0=1 kvsatdpl=0                   wdpl=0 kvth0dpl_b1=-0.000            kvth0dpl_b2=-0.000            dplbinflg=0 ku0dpl_b1=0                 ku0dpl_b2=0 keta0dpl_b1=0                  keta0dpl_b2=0 kvth0dpx=0                  wkvth0dpx=0e-07               wdpxkvth0=1 lkvth0dpx=0.0e-8              ldpxkvth0=1.0                 pkvth0dpx=0.0e-18 ku0dpx=0                   wku0dpx=0e-9                wdpxku0=1 lku0dpx=0e-8                ldpxku0=1.0                 pku0dpx=0.0e-18 keta0dpx=0.00                wketa0dpx=0e-7                wdpxketa0=1 kvsatdpx=0.00                wdpx=0 kvth0dpx_b1=-0.000            kvth0dpx_b2=-0.000            dpxbinflg=0 ku0dpx_b1=0                 ku0dpx_b2=0 keta0dpx_b1=0                  keta0dpx_b2=0 kvth0dps=0                   wkvth0dps=0                   wdpskvth0=1 lkvth0dps=-0.0e-9             ldpskvth0=1.0                 pkvth0dps=0 ku0dps=0                   wku0dps=-0.0e-9             wdpsku0=1 lku0dps=0e-15               ldpsku0=2.0                 pku0dps=0e-23 keta0dps=0                   wketa0dps=0                   wdpsketa0=1 kvsatdps=0                   wdps=0 kvth0dps_b1=-0.000            kvth0dps_b2=-0.000            dpsbinflg=0 ku0dps_b1=0                 ku0dps_b2=0 keta0dps_b1=0                  keta0dps_b2=0 kvth0dpa=-0.007              wkvth0dpa=-0.0e-10            wdpakvth0=1 lkvth0dpa=-1e-8               ldpakvth0=1.0                 pkvth0dpa=0.0e-19 ku0dpa=-0.02               wku0dpa=2e-9                wdpaku0=1 lku0dpa=-4.0e-8             ldpaku0=1.0                 pku0dpa=-0.0e-18 keta0dpa=0.00                wketa0dpa=0e-7                wdpaketa0=1 ka0dpa=0.0                 wka0dpa=0                   wdpaka0=1 lka0dpa=0.0e-7              ldpaka0=1.0                 pka0dpa=0.0e-14 kvsatdpa=0                   wdpa=0 kvth0dpa_b1=0.006             kvth0dpa_b2=-0.006            dpabinflg=0 ku0dpa_b1=-0.04             ku0dpa_b2=0.04 keta0dpa_b1=0                  keta0dpa_b2=0 ka0dpa_b1=0                 ka0dpa_b2=0 spbref=5.31e-7             spbmax='1.6e-6+1.2e-6+0.2e-6'    spbmin='1.98e-7+1.98e-7+0.2e-6' pse_mode=1 kvth0dp2=0                   wkvth0dp2=-0.0e-8             wdp2kvth0=1 lkvth0dp2=0e-9                ldp2kvth0=1.0                 pkvth0dp2=0.0e-19 ku0dp2=0.0                 wku0dp2=-0.0e-8             wdp2ku0=1 lku0dp2=0e-5                ldp2ku0=0.5                 pku0dp2=0 keta0dp2=0.00                wketa0dp2=-0e-9               wdp2keta0=1 kvsatdp2=0                   wdp2=0 kvth0dp2l=-0.00              wkvth0dp2l=-0.0e-8            wdp2lkvth0=1 lkvth0dp2l=0.0e-9             ldp2lkvth0=1                  pkvth0dp2l=0 ku0dp2l=0.00               wku0dp2l=-0.0e-8            wdp2lku0=1 lku0dp2l=0.0e-9             ldp2lku0=1.0                pku0dp2l=0 keta0dp2l=0.00               wketa0dp2l=-0e-9              wdp2lketa0=1 kvsatdp2l=0                  wdp2l=0 kvth0dp2l_b1=0.016            kvth0dp2l_b2=-0.016           dp2lbinflg=0 ku0dp2l_b1=-0.04            ku0dp2l_b2=0.04 keta0dp2l_b1=0                 keta0dp2l_b2=0 kvth0dp2a=0.00               wkvth0dp2a=-0.0e-9            wdp2akvth0=1 lkvth0dp2a=0.0e-9             ldp2akvth0=1.0                pkvth0dp2a=-0.0e-17 ku0dp2a=0.00               wku0dp2a=0e-9               wdp2aku0=1 lku0dp2a=0.0e-5             ldp2aku0=0.5                pku0dp2a=-0.0e-18 keta0dp2a=0.00               wketa0dp2a=0e-7               wdp2aketa0=1 ka0dp2a=0                  wka0dp2a=0                  wdp2aka0=1 lka0dp2a=0                  ldp2aka0=1.0                pka0dp2a=0.0e-14 kvsatdp2a=0.00               wdp2a=0 kvth0dp2a_b1=-0.000           kvth0dp2a_b2=-0.000           dp2abinflg=0 ku0dp2a_b1=0                ku0dp2a_b2=0 keta0dp2a_b1=0                 keta0dp2a_b2=0 ka0dp2a_b1=0                 ka0dp2a_b2=0 enxref=1.0e-5              enxmax=1.0e-5              enxmin=1e-6 kvth0enx=0           	 wkvth0enx=0                   wenxkvth0=1 lkvth0enx=0          	 lenxkvth0=1                   pkvth0enx=0 ku0enx=0         		 wku0enx=0      		 wenxku0=1 lku0enx=0          	 lenxku0=1                   pku0enx=0 keta0enx=0                   wketa0enx=0                   wenxketa0=1 ka0enx=0                   wka0enx=0                   wenxka0=1 lka0enx=0          	 lenxka0=1                   pka0enx=0 kvsatenx=0                   wenx=0                   ku0enx0=0 eny0=2.0e-6 enyref=2.0e-6              enymax=2.0e-6              enymin=0.05e-6 kvth0eny=0          	 wkvth0eny=0       		 wenykvth0=1 lkvth0eny=0        		 lenykvth0=1                   pkvth0eny=0 ku0eny=0          	 wku0eny=0        		 wenyku0=1 ku0eny0=0          	 wku0eny0=0                   weny0ku0=1 lku0eny=0       		 lenyku0=1                 	 pku0eny=0 keta0eny=0               	 wketa0eny=0                   wenyketa0=1 ka0eny=0              	 wka0eny=0             	 wenyka0=1 lka0eny=0      		 lenyka0=1                	 pka0eny=0 kvsateny=0               	 weny=0 kvth0eny1=0             	 wkvth0eny1=0        		 weny1kvth0=1 lkvth0eny1=0             	 leny1kvth0=1                  pkvth0eny1=0 ku0eny1=0        		 wku0eny1=0            	 weny1ku0=1 lku0eny1=0      		 leny1ku0=1                	 pku0eny1=0 keta0eny1=0              	 wketa0eny1=0                  weny1keta0=1 ka0eny1=0                  wka0eny1=0                  weny1ka0=1 lka0eny1=0                  leny1ka0=1                	 pka0eny1=0 kvsateny1=0               	 weny1=0 rx_mode=0 rxref=1.8126e-5           ringxmax=0.8126e-5           ringxmin=0 kvth0rx=0              	 wkvth0rx=0          	 wrxkvth0=1 lkvth0rx=0              	 lrxkvth0=1                	 pkvth0rx=0 ku0rx=0              	 wku0rx=0           	 wrxku0=1 lku0rx=0        		 lrxku0=1                   pku0rx=0 keta0rx=0                	 wketa0rx=0                   wrxketa0=1 kvsatrx=0                	 wrx=0                   ku0rx0=0 ry_mode=0 ryref=1.8027e-5           ringymax=1.6027e-5           ringymin=0 kvth0ry=0           	 wkvth0ry=0           	 wrykvth0=1 lkvth0ry=0              	 lrykvth0=1                 	 pkvth0ry=0 ku0ry=0          	 wku0ry=0           	 wryku0=1 lku0ry=0        		 lryku0=1                 	 pku0ry=0 keta0ry=0                	 wketa0ry=0                   wryketa0=1 kvsatry=0                   wry=0 kvth0ry0=0                	 ku0ry0=0 sfxref=8.26e-7           sfxmax=3e-6               minwodx=0.53e-6 sfxmin=0.189e-6 lrefodx=5e-8              lodxref=1                 wodx=1e-6 kvth0odxa=-0.200            lkvth0odxa=1.0e-13           lodxakvth0=2.0 wkvth0odxa=5.0e-12           wodxakvth0=2.0               pkvth0odxa=0.0e-16 ku0odxa=-1.20             lku0odxa=2.0e-13           lodxaku0=2.0 wku0odxa=5.0e-12           wodxaku0=1.0               pku0odxa=0.0e-16 keta0odx=0.0               wketa0odx=0                 wodxketa0=1 kvsatodx=0.0 kvth0odxb=-0.00             lkvth0odxb=-0.0e-7           lodxbkvth0=0.5 wkvth0odxb=-0.0e-5           wodxbkvth0=1.0               pkvth0odxb=0.0e-16 ku0odxb=-0.00             lku0odxb=0.0e-7            lodxbku0=0.5 wku0odxb=-0.0e-5           wodxbku0=1.0               pku0odxb=0.0e-16 lrefodx1=5e-8              lodx1ref=1                 r_sodx1=1 kvth0odx1a=-0.000            lkvth0odx1a=1.0e-13           lodx1akvth0=2.0 wkvth0odx1a=0.0e-7            wodx1akvth0=1.0               pkvth0odx1a=0.0e-16 ku0odx1a=-0.00             lku0odx1a=1.0e-13           lodx1aku0=2.0 wku0odx1a=0.0e-7            wodx1aku0=1.0               pku0odx1a=0.0e-16 keta0odx1=0.00              wketa0odx1=0                 wodx1keta0=1 kvsatodx1=0.0 kvth0odx1b=-0.0005           lkvth0odx1b=0.0e-7            lodx1bkvth0=0.5 wkvth0odx1b=-2.0e-15          wodx1bkvth0=2.0               pkvth0odx1b=0.0e-16 ku0odx1b=-0.00             lku0odx1b=0.0e-7            lodx1bku0=0.5 wku0odx1b=-1.5e-14          wodx1bku0=2.0               pku0odx1b=0.0e-16 sfyref=7.9e-7 sfymin=0.15e-6 sfymax=3e-6              minwody=0e-7              wody=1e-6 kvth0odya=-0.000            lkvth0odya=1.0e-13           lodyakvth0=2.0 wkvth0odya=0.0e-6            wodyakvth0=1.0               pkvth0odya=0.0e-16 ku0odya=-2.00             lku0odya=2.0e-13           lodyaku0=2.0 wku0odya=0.0e-6            wodyaku0=1.0               pku0odya=0.0e-16 keta0ody=0.00              wketa0ody=0                 wodyketa0=1 kvsatody=0.0 lrefody=5e-8              lodyref=1 kvth0odyb=-0.00             lkvth0odyb=-3.0e-9           lodybkvth0=1.0 wkvth0odyb=-7.0e-8           wodybkvth0=1.0               pkvth0odyb=0.0e-15 ku0odyb=0.10              lku0odyb=0.0e-9            lodybku0=0.8 wku0odyb=-0.0e-5           wodybku0=1.0               pku0odyb=0.0e-13 web_mac=-0  wec_mac=-0 kvsatwe=-0 lodflag=1    pseflag=1 ceslflag=0 oseflag=1 wpeflag=0 )
.model nch_na18ud15_mac.1 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=9e-006                     wmax=0.00090001                 vth0=-0.1312 k2=0.0147                     minv=-0.21803                   cit=0.0001 voff=-0.118                     eta0=0.12                       etab=0.01 u0=0.042179                   ua=-3e-011                    ub=2.78e-018 uc=6.5485e-011                vsat=80000                      a0=6.7 ags=1.15                       keta=-0.028                     pclm=1 pdiblc2=0.0021                     tvoff=0.001824                   ltvoff=0 wtvoff=0                          ptvoff=0                          kt1=-0.17 kt2=-0.0024                    ute=-1.86                      ua1=8e-010 ub1=-2.6182e-018               uc1=-7.1e-011                  at=80000 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=0                          wk2=0 wvoff=0                          weta0=0                          wu0=0 wa0=0                          wags=0                          wpdiblc2=0 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wvsat=0                          pvsat=0 wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18ud15_mac.2 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.13125028 k2=0.016409444                minv=-0.21803                   cit=0.0001 voff=-0.122525                  eta0=0.11698333                 etab=0.01 u0=0.041860993                ua=-3.2513889e-011            ub=2.7875417e-018 uc=7.2587842e-011             vsat=80000                      a0=7.0066944 ags=1.0557292                  keta=-0.024983333               pclm=0.84916667 pdiblc2=0.0013709722               tvoff=0.00145446                 ltvoff=3.32957e-009 wtvoff=0                          ptvoff=0                          kt1=-0.16874306 kt2=0.000274275                ute=-1.858014                  ua1=7.8464014e-010 ub1=-2.3012388e-018            uc1=-7.5005429e-011            at=80502.778 lvth0=4.5300278e-010             lk2=-1.5402094e-008            lvoff=4.077025e-008 leta0=2.7180167e-008             lu0=2.8652426e-009             lua=2.2650139e-017 lub=-6.7950417e-026            luc=-6.3996608e-017            la0=-2.7633169e-006 lags=8.4938021e-007             lketa=-2.7180167e-008            lpclm=1.3590083e-006 lpdiblc2=6.5685403e-009             lkt1=-1.1325069e-008            lkt2=-2.4095218e-008 lute=-1.789361e-008             lua1=1.3839235e-016             lub1=-2.8558201e-024 luc1=3.6088919e-017             lat=-0.0045300278              lvsat=0 lcit=0                          wvth0=0                          wk2=0 wvoff=0                          weta0=0                          wu0=0 wa0=0                          wags=0                          wpdiblc2=0 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wvsat=0                          pvsat=0 wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18ud15_mac.3 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.13069722 k2=0.0060833333               minv=-0.21803                   cit=0.0001 voff=-0.1                       eta0=0.19558333                 etab=0.0061865139 u0=0.043737694                ua=-4.8611111e-012            ub=2.9392361e-018 uc=4.3058467e-011             vsat=78788.889                  a0=6.0552778 ags=1.7142361                  keta=-0.018805556               pclm=1.7513889 pdiblc2=0.0072708333               tvoff=0.00142102                 ltvoff=3.3901e-009 wtvoff=0                          ptvoff=0                          kt1=-0.18256944 kt2=-0.025206639               ute=-2.034125                  ua1=5.0579028e-010 ub1=-4.0326089e-018            uc1=-2.5047216e-011            at=149092.22 lvth0=-5.4802778e-010            lk2=3.2881667e-009             lvoff=0 leta0=-1.1508583e-007            lu0=-5.3158694e-010            lua=-2.7401389e-017 lub=-3.4251736e-025            luc=-1.0548439e-017            la0=-1.0412528e-006 lags=-3.4251736e-007            lketa=-3.8361944e-008            lpclm=-2.7401389e-007 lpdiblc2=-4.1102083e-009            lkt1=1.3700694e-008             lkt2=2.2025236e-008 lute=3.0086725e-007             lua1=6.431106e-016              lub1=2.7795969e-025 luc1=-5.4335447e-017            lat=-0.12867692                letab=6.9024099e-009 lvsat=0.0021921111               lcit=0                          wvth0=0 wk2=0                          wvoff=0                          weta0=0 wu0=0                          wa0=0                          wags=0 wpdiblc2=0                          pvth0=0                          pk2=0 pvoff=0                          peta0=0                          pu0=0 pags=0                          ppdiblc2=0                          wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18ud15_mac.4 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=9e-006                     wmax=0.00090001                 vth0=-0.13870278 k2=0.012547222                minv=-0.51426806                cit=-0.0012789294 voff=-0.089861111               eta0=0.15083333                 etab=0.017626972 u0=0.041222222                ua=-3e-011                    ub=2.8277778e-018 uc=4.6510861e-011             vsat=81083.889                  a0=4.8972222 ags=1.9069444                  keta=-0.082388889               pclm=1.9055556 pdiblc2=0.0075555556               tvoff=-0.000205283               ltvoff=5.16277e-009 wtvoff=0                          ptvoff=0                          kt1=-0.18778361 kt2=0.01633425                 ute=-1.7603306                 ua1=1.5728347e-009 ub1=-5.3544e-018               uc1=-2.0737209e-010            at=83202.758 lvth0=8.1780278e-009             lk2=-3.7574722e-009            lvoff=-1.1051389e-008 leta0=-6.6308333e-008            lu0=2.2102778e-009             lub=-2.2102778e-025 luc=-1.4311549e-017            la0=2.2102778e-007             lags=-5.5256944e-007 lketa=3.0943889e-008             lpclm=-4.4205556e-007            lpdiblc2=-4.4205556e-009 lkt1=1.9384136e-008             lkt2=-2.3254333e-008            lute=2.4313056e-009 lua1=-5.1996785e-016            lub1=1.718712e-024              luc1=1.4439866e-016 lat=-0.056857407               letab=-5.5676897e-009            lvsat=-0.00030943889 lminv=3.2289948e-007             lcit=1.5030331e-009             wvth0=0 wk2=0                          wvoff=0                          weta0=0 wu0=0                          wa0=0                          wags=0 wpdiblc2=0                          pvth0=0                          pk2=0 pvoff=0                          peta0=0                          pu0=0 pags=0                          ppdiblc2=0                          wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=0 tmimodel=1 )
.model nch_na18ud15_mac.5 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.131375 k2=0.016125                   minv=-0.1725375                 cit=0.0001 voff=-0.123                     eta0=0.13312675                 etab=0.01 u0=0.04247375                 ua=-3.8e-011                  ub=2.8375e-018 uc=7.152075e-011              vsat=80000                      a0=7.0225 ags=1.1325                     keta=-0.031875                  pclm=1 pdiblc2=0.002125                   tvoff=0.00123                    ltvoff=0 wtvoff=5.346e-009                 ptvoff=0                          kt1=-0.17125 kt2=0.00088025                 ute=-1.865                     ua1=7.6451e-010 ub1=-2.50685e-018              uc1=-8.20675e-011              at=82500 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=1.575e-009                 wk2=-1.2825e-008 wminv=-4.094325e-007             wvoff=4.5e-008                   weta0=-1.1814075e-007 wu0=-2.65275e-009              wua=7.2e-017                   wub=-5.175e-025 wuc=-5.432175e-017             wa0=-2.9025e-006               wags=1.575e-007 wketa=3.4875e-008                wpdiblc2=-2.25e-010                 wkt1=1.125e-008 wkt2=-2.952225e-008             wute=4.5e-008                   wua1=3.1941e-016 wub1=-1.00215e-024              wuc1=9.96075e-017               wat=-0.0225 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wvsat=0                          pvsat=0 wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.6 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.13102934 k2=0.018431493                minv=-0.17283225                cit=0.0001 voff=-0.12909618                eta0=0.13099441                 etab=0.01 u0=0.042246432                ua=-3.9382639e-011            ub=2.8506979e-018 uc=8.090697e-011              vsat=80000                      a0=7.2999705 ags=1.0385434                  keta=-0.030460937               pclm=0.84288194 pdiblc2=0.0015279514               tvoff=0.00072232                 ltvoff=4.5742e-009 wtvoff=6.58924e-009               ptvoff=-1.12016e-014              kt1=-0.16999306 kt2=0.0047345602               ute=-1.8608018                 ua1=7.3182065e-010 ub1=-2.1329907e-018            uc1=-9.0283299e-011            at=83243.734 lvth0=-3.1143941e-009            lk2=-2.0781502e-008            lvoff=5.4926587e-008 leta0=1.9212414e-008             lu0=2.0481388e-009             lua=1.2457576e-017 lub=-1.1891323e-025            luc=-8.4569843e-017            la0=-2.5000091e-006 lags=8.4654894e-007             lketa=-1.2740703e-008            lpclm=1.4156337e-006 lpdiblc2=5.379408e-009              lkt1=-1.1325069e-008            lkt2=-3.4727335e-008 lute=-3.7825732e-008            lua1=2.9453108e-016             lub1=-3.368472e-024 luc1=7.4024346e-017             lat=-0.0067010436              lvsat=0 lminv=2.6557288e-009             lcit=0                          wvth0=-1.9884375e-009 wk2=-1.8198438e-008            wminv=-4.0677972e-007            wvoff=5.9140625e-008 weta0=-1.2609966e-007            wu0=-3.4689469e-009            wua=6.181875e-017 wub=-5.6840625e-025            wuc=-7.4872151e-017            wa0=-2.6394844e-006 wags=1.5467187e-007             wketa=4.9298438e-008             wpdiblc2=-1.4128125e-009 wkt1=1.125e-008                 wkt2=-4.0142566e-008            wute=2.509e-008 wua1=4.7537544e-016             wub1=-1.5142329e-024            wuc1=1.3750082e-016 wat=-0.024668606               pvth0=3.2106572e-014             pk2=4.8414672e-014 pminv=-2.3901559e-014            pvoff=-1.2740703e-013            peta0=7.1709773e-014 pu0=7.3539338e-015             pua=9.1733062e-023             pub=4.5866531e-031 puc=1.8515911e-022             pa0=-2.3697708e-012            pags=2.5481406e-014 pketa=-1.2995517e-013            wpclm=5.65625e-008               ppclm=-5.0962812e-013 ppdiblc2=1.0702191e-014             pkt1=-5.4065258e-028            pkt2=9.5689051e-014 pute=1.793891e-013              pua1=-1.4052486e-021            pub1=4.6138673e-030 puc1=-3.4141884e-022            pat=1.9539142e-008             wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.7 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.13199306 k2=0.0034018229               minv=-0.171365                  cit=0.0001 voff=-0.098606181               eta0=0.21595457                 etab=0.013821434 u0=0.044075903                ua=-1.3576389e-011            ub=3.0026215e-018 uc=3.5714311e-011             vsat=78486.111                  a0=6.9122396 ags=1.6671007                  keta=-0.015548611               pclm=1.8142361 pdiblc2=0.0066194444               tvoff=0.00130567                 ltvoff=3.51834e-009 wtvoff=1.03815e-009               ptvoff=-1.15415e-015              kt1=-0.18646875 kt2=-0.032801376               ute=-2.0482278                 ua1=5.4561632e-010 ub1=-4.1522642e-018            uc1=2.7273593e-012             at=153084.33 lvth0=-1.3700694e-009            lk2=6.4222005e-009             lvoff=-2.6031319e-010 leta0=-1.3456548e-007            lu0=-1.263204e-009             lua=-3.4251736e-017 lub=-3.9389496e-025            luc=-2.7711299e-018            la0=-1.7982161e-006 lags=-2.9113976e-007            lketa=-3.9732014e-008            lpclm=-3.4251736e-007 lpdiblc2=-3.8361944e-009            lkt1=1.8495937e-008             lkt2=3.321271e-008 lute=3.0141528e-007             lua1=6.3156091e-016             lub1=2.8641302e-025 luc1=-9.4324945e-017            lat=-0.13311252                letab=-6.9167956e-009 lvsat=0.0027401389               lcit=0                          wvth0=1.16625e-008 wk2=2.4133594e-008             wminv=-4.19985e-007              wvoff=-1.2544375e-008 weta0=-1.8334112e-007            wu0=-3.043875e-009             wua=7.84375e-017 wub=-5.7046875e-025            wuc=6.6097401e-017             wa0=-7.7126563e-006 wags=4.2421875e-007             wketa=-2.93125e-008              wpdiblc2=5.8625e-009 wkt1=3.509375e-008              wkt2=6.8352633e-008             wute=1.26925e-007 wua1=-3.5843437e-016            wub1=1.0768981e-024             wuc1=-2.4997118e-016 wat=-0.035928969               pvth0=7.398375e-015              pk2=-2.8206305e-014 pvoff=2.3428188e-015             peta0=1.7531683e-013             pu0=6.5845538e-015 pua=6.1653125e-023             pub=4.6239844e-031             puc=-6.9995779e-023 pa0=6.8126703e-012             pags=-4.6239844e-013            pketa=1.2330625e-014 wpclm=-5.65625e-007              ppclm=6.1653125e-013             ppdiblc2=-2.466125e-015 pkt1=-4.3157188e-014            pkt2=-1.0068726e-013            pute=-4.93225e-015 pua1=1.0394717e-022             pub1=-7.6079956e-032            puc1=3.5990548e-022 pat=3.9920398e-008             wetab=-6.8714281e-008            petab=1.2437285e-013 wvsat=0.002725                   pvsat=-4.93225e-009              wcit=0 pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.8 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=1.8e-006                   wmax=9e-006                     vth0=-0.14288194 k2=0.016915964                minv=-0.44702111                cit=-0.0010545153 voff=-0.10410708                eta0=0.1609375                  etab=0.0023880556 u0=0.040239319                ua=-4.6776333e-011            ub=2.7755903e-018 uc=6.2007061e-011             vsat=81599.208                  a0=3.9190972 ags=1.9829861                  keta=-0.08636475                pclm=1.8548611 pdiblc2=0.0068006944               tvoff=-0.00114478                ltvoff=6.18933e-009 wtvoff=8.45551e-009               ptvoff=-9.23907e-015              kt1=-0.20338924 kt2=0.024415389                ute=-1.8393771                 ua1=1.5108502e-009 ub1=-5.6653264e-018            uc1=-2.6200832e-010            at=87361.08 lvth0=1.0498819e-008             lk2=-8.3082131e-009            lvoff=5.7356708e-009 leta0=-7.4596875e-008            lu0=2.9186718e-009             lua=1.9362033e-018 lub=-1.464309e-025             luc=-3.1430227e-017            la0=1.464309e-006 lags=-6.3545486e-007            lketa=3.7457578e-008             lpclm=-3.8679861e-007 lpdiblc2=-4.0337569e-009            lkt1=3.6939267e-008             lkt2=-2.9153564e-008 lute=7.3768021e-008             lua1=-4.2054403e-016            lub1=1.9356508e-024 luc1=1.9423695e-016             lat=-0.06147418                letab=5.5455869e-009 lvsat=-0.00065313708             lminv=3.0046516e-007             lcit=1.2584216e-009 wvth0=3.76125e-008               wk2=-3.9318675e-008            wminv=-6.052225e-007 wvoff=1.2821375e-007             weta0=-9.09375e-008              wu0=8.846125e-009 wua=1.50987e-016               wub=4.696875e-025              wuc=-1.394658e-016 wa0=8.803125e-006              wags=-6.84375e-007              wketa=3.578275e-008 wpdiblc2=6.79375e-009               wkt1=1.4045062e-007             wkt2=-7.273025e-008 wute=7.1141875e-007             wua1=5.5786062e-016             wub1=2.7983375e-024 wuc1=4.9172609e-016             wat=-0.037424894               pvth0=-2.0887125e-014 pk2=4.0956668e-014             pminv=2.0190888e-013             pvoff=-1.5108354e-013 peta0=7.4596875e-014             pu0=-6.3755462e-015            pua=-1.742583e-023 pub=-6.7137188e-031            puc=1.5406811e-022             pa0=-1.1189531e-011 pags=7.4596875e-013             pketa=-5.8623197e-014            wpclm=4.5625e-007 ppclm=-4.973125e-013             ppdiblc2=-3.4811875e-015            pkt1=-1.5799618e-013 pkt2=5.3093083e-014             pute=-6.4203044e-013            pua1=-8.9481438e-022 pub1=-1.9524489e-030            puc1=-4.4854454e-022            pat=4.1550957e-008 wetab=1.3715025e-007             petab=-1.0001949e-013            wvsat=-0.004637875 pvsat=3.0932837e-009             wcit=-2.0197275e-009            pcit=2.201503e-015 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.9 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.1233 k2=0.0075                     minv=-0.28585                   cit=0.0001 voff=-0.098363                  eta0=0.067493                   etab=0.01 u0=0.03995                    ua=3.5e-013                   ub=2.49e-018 uc=5.3288e-011                vsat=80000                      a0=4.525 ags=1.52                       keta=-0.00425                   pclm=1 pdiblc2=0.00185                    tvoff=0.004425                   ltvoff=0 wtvoff=-4.05e-010                 ptvoff=0                          kt1=-0.1725 kt2=-0.015521                  ute=-1.975                     ua1=5.327e-010 ub1=-2.709e-018                uc1=-5.478e-012                at=62500 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=-1.296e-008                wk2=2.7e-009 wminv=-2.0547e-007               wvoff=6.534e-010                 weta0=0 wu0=1.89e-009                  wua=2.97e-018                  wub=1.08e-025 wuc=-2.15028e-017              wa0=1.593e-006                 wags=-5.4e-007 wketa=-1.485e-008                wpdiblc2=2.7e-010                   wkt1=1.35e-008 wute=2.43e-007                  wua1=7.36668e-016               wub1=-6.3828e-025 wuc1=-3.82536e-017              wat=0.0135                     pvth0=0 pk2=0                          pvoff=0                          peta0=0 pu0=0                          pags=0                          ppdiblc2=0 wvsat=0                          pvsat=0                          wcit=0 pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.10 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.12478319 k2=0.006934375                minv=-0.28290246                cit=0.0001 voff=-0.098865778               eta0=0.081639407                etab=0.058360938 u0=0.038595768                ua=-7.1036806e-012            ub=2.4145833e-018 uc=5.4861192e-011             vsat=80000                      a0=4.5988832 ags=1.4659514                  keta=0.00366875                 pclm=0.98743056 pdiblc2=-0.00050048611             tvoff=0.00514498                 ltvoff=-6.487e-009 wtvoff=-1.37154e-009              ptvoff=8.70853e-015               kt1=-0.17312847 kt2=-0.020635664               ute=-1.9741704                 ua1=6.0054986e-010 ub1=-2.5752485e-018            uc1=2.6196573e-011             at=60098.105 lvth0=1.3363582e-008             lk2=5.0962812e-009             lvoff=4.5300278e-009 leta0=-1.2745913e-007            lu0=1.220163e-008              lua=6.7157662e-017 lub=6.7950417e-025             luc=-1.4174457e-017            la0=-6.6568758e-007 lags=4.8697799e-007             lketa=-7.1347937e-008            lpclm=1.1325069e-007 lpdiblc2=2.117788e-008              lkt1=5.6625347e-009             lkt2=4.6083123e-008 lute=-7.4745458e-009            lua1=-6.1132725e-016            lub1=-1.2051006e-024 luc1=-2.853879e-016             lat=0.021641075                letab=-4.3573205e-007 lvsat=0                          lminv=-2.6557288e-008            lcit=0 wvth0=-1.32315e-008              wk2=2.496375e-009              wminv=-2.0865334e-007 wvoff=4.7259e-009                weta0=-3.726066e-008             wu0=3.1022475e-009 wua=3.716625e-018              wub=2.166e-025                 wuc=-2.7989749e-017 wa0=2.2224727e-006             wags=-6.146625e-007             wketa=-1.2135e-008 wpdiblc2=2.238375e-009              wkt1=1.689375e-008              wkt2=5.5238372e-009 wute=2.291535e-007              wua1=7.1166285e-016             wub1=-7.1816887e-025 wuc1=-7.2162945e-017            wat=0.016993526                pvth0=2.446215e-015 pk2=1.8346612e-015             pminv=2.8681871e-014             pvoff=-3.6693225e-014 peta0=3.3571855e-013             pu0=-1.092235e-014             pua=-6.7270913e-024 pub=-9.78486e-031              puc=5.8447415e-023             pa0=-5.6715495e-012 pags=6.7270913e-013             pketa=-2.446215e-014             wpclm=-2.03625e-007 ppclm=1.8346612e-012             ppdiblc2=-1.7735059e-014            pkt1=-3.0577687e-014 pkt2=-4.9769773e-014            pute=1.2475697e-013             pua1=2.252964e-022 pub1=7.1979876e-031             puc1=3.055232e-022              pat=-3.1476671e-008 wetab=-8.7049687e-008            petab=7.8431768e-013             wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.11 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.10778681 k2=0.0077630208               minv=-0.297575                  cit=0.0011922708 voff=-0.079389278               eta0=-0.024780278               etab=-0.49136729 u0=0.043963903                ua=3e-011                     ub=2.7748611e-018 uc=4.7788307e-011             vsat=80000                      a0=2.4236681 ags=2.1967361                  keta=0.00171875                 pclm=-0.76666667 pdiblc2=0.018618056                tvoff=-0.00283102                ltvoff=7.94955e-009 wtvoff=8.48418e-009               ptvoff=-9.13033e-015              kt1=-0.18968056 kt2=0.036212273                ute=-2.4344347                 ua1=-1.1502866e-009 ub1=-2.5159729e-018            uc1=-2.4003129e-010            at=136366.77 lvth0=-1.7399882e-008            lk2=3.5964323e-009             lvoff=-3.0722437e-008 leta0=6.5160503e-008             lu0=2.485306e-009              lub=2.7401389e-026 luc=-1.3725356e-018            la0=3.2714518e-006             lags=-8.3574236e-007 lketa=-6.7818438e-008            lpclm=3.2881667e-006             lpdiblc2=-1.3426681e-008 lkt1=3.5621806e-008             lkt2=-5.6811642e-008            lute=8.2560385e-007 lua1=2.5576867e-015             lub1=-1.3123895e-024            luc1=1.9648454e-016 lat=-0.11640521                letab=5.5927605e-007             lvsat=0 lcit=-1.9770102e-009            wvth0=-3.190875e-008             wk2=1.6283437e-008 wminv=-1.92807e-007              wvoff=-4.71348e-008              weta0=2.499816e-007 wu0=-2.842275e-009             wub=-1.605e-025                wuc=4.4364208e-017 wa0=3.667725e-007              wags=-5.29125e-007              wketa=-6.039375e-008 wpdiblc2=-1.5735e-008               wkt1=4.0875e-008                wkt2=-5.5871934e-008 wute=8.220975e-007              wua1=2.6941909e-015             wub1=-1.8684263e-024 wuc1=1.869944e-016              wat=-0.0058373625              pvth0=3.6252037e-014 pk2=-2.3119922e-014            pvoff=5.7174642e-014             peta0=-1.8418994e-013 pu0=-1.6276425e-016            pub=-2.95935e-031              puc=-7.2513249e-023 pa0=-2.312732e-012             pags=5.1788625e-013             pketa=6.2886187e-014 wpclm=4.08e-006                  ppclm=-5.9187e-012               ppdiblc2=1.479675e-014 pkt1=-7.398375e-014             pkt2=6.1356573e-014             pute=-9.4847168e-013 pua1=-3.3630793e-021            pub1=2.8017646e-030             puc1=-1.6355159e-022 pat=9.8472371e-009             wetab=8.4062543e-007             petab=-8.9477427e-013 wvsat=0                          pvsat=0                          wcit=-1.9660875e-009 pcit=3.5586184e-015 lmin_flag=1                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.12 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=1.08e-006                  wmax=1.8e-006                   vth0=-0.13246944 k2=0.011388972                minv=-0.40418542                cit=-0.0043611278 voff=-0.072240972               eta0=-0.0045416667              etab=0.067924806 u0=0.050033917                ua=4.7763333e-011             ub=3.5806944e-018 uc=-1.6496971e-011            vsat=79022.611                  a0=11.457639 ags=1.1765278                  keta=-0.11733861                pclm=3.7708333 pdiblc2=0.00995                    tvoff=0.00489234                 ltvoff=-4.6891e-010 wtvoff=-2.41132e-009              ptvoff=2.74576e-015               kt1=-0.087548611 kt2=-0.11938245                ute=-1.0819486                 ua1=2.9816632e-009 ub1=-4.7592361e-018            uc1=2.6294189e-010             at=62357.097 lvth0=9.5041944e-009             lk2=-3.5585472e-010            lvoff=-3.851409e-008 leta0=4.3100417e-008             lu0=-4.1310092e-009            lua=-1.9362033e-017 lub=-8.5095694e-025            luc=6.8698417e-017             la0=-6.5755764e-006 lags=2.7628472e-007             lketa=6.1954086e-008             lpclm=-1.6577083e-006 lpdiblc2=-3.9785e-009               lkt1=-7.5702014e-008            lkt2=1.1278661e-007 lute=-6.4860601e-007            lua1=-1.9461385e-015            lub1=1.1327674e-024 luc1=-3.5175624e-016            lat=-0.035734666               letab=-5.0352338e-008 lvsat=0.0010653539               lminv=1.1620535e-007             lcit=4.0761943e-009 wvth0=1.887e-008                 wk2=-2.937009e-008             wminv=-6.8232675e-007 wvoff=7.085475e-008              weta0=2.06925e-007               wu0=-8.78415e-009 wua=-1.91844e-017              wub=-9.795e-025                wuc=1.8414585e-018 wa0=-4.76625e-006              wags=7.6725e-007                wketa=9.15357e-008 wpdiblc2=1.125e-009                 wkt1=-6.80625e-008              wkt2=1.8610586e-007 wute=-6.519525e-007             wua1=-2.0896027e-015            wub1=1.167375e-024 wuc1=-4.5318429e-016            wat=0.007582275                pvth0=-1.90968e-014 pk2=2.6642423e-014             pminv=5.3357653e-013             pvoff=-7.1433968e-014 peta0=-1.3725825e-013            pu0=6.3138795e-015             pua=2.0910996e-023 pub=5.96775e-031               puc=-2.6163452e-023            pa0=3.2822625e-012 pags=-8.951625e-013             pketa=-1.0271691e-013            wpclm=-2.9925e-006 ppclm=1.790325e-012              ppdiblc2=-3.58065e-015              pkt1=4.4758125e-014 pkt2=-2.0239923e-013            pute=6.5824283e-013             pua1=1.8512557e-021 pub1=-5.0725875e-031            puc1=5.3424318e-022             pat=-4.7801678e-009 wetab=1.91841e-008               petab=5.96775e-016               wvsat=0 pvsat=0                          wcit=3.932175e-009              pcit=-2.8704878e-015 lmin_flag=0                          lmax_flag=1                          wmin_flag=1 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.13 nmos ( level=54                         lmin=9e-006                     lmax=0.00090001 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.14033571 k2=0.012766429                minv=-0.4761                    cit=0.0001 voff=-0.096329429               eta0=0.067493                   etab=0.013051357 u0=0.041477857                ua=-1.5145e-011               ub=2.7757143e-018 uc=2.1125857e-011             vsat=80000                      a0=7.2857143 ags=1.0574286                  keta=-0.024964286               pclm=1 pdiblc2=0.0021714286               tvoff=0.00405286                 ltvoff=0 wtvoff=-3.08571e-012              ptvoff=0                          kt1=-0.13682143 kt2=-0.015521                  ute=-1.7142857                 ua1=1.5591571e-009 ub1=-3.8617143e-018            uc1=-3.8385143e-011            at=75000 lvth0=0                          lk2=0                          lvoff=0 leta0=0                          lu0=0                          luc=0 la0=0                          lags=0                          lketa=0 lpdiblc2=0                          lkt2=0                          lvsat=0 lcit=0                          wvth0=5.4385714e-009             wk2=-2.9877429e-009 wvoff=-1.5428571e-009            weta0=0                          wu0=2.3991429e-010 wua=1.97046e-017               wub=-2.0057143e-025            wuc=1.3232314e-017 wa0=-1.3885714e-006            wags=-4.0422857e-008            wketa=7.5214286e-009 wpdiblc2=-7.7142857e-011            wkt1=-2.5032857e-008            wute=-3.8571429e-008 wua1=-3.7190571e-016            wub1=6.0665143e-025             wuc1=-2.7138857e-018 pvth0=0                          pk2=0                          pvoff=0 peta0=0                          pu0=0                          pags=0 ppdiblc2=0                          wetab=-3.2954657e-009            wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=0                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.14 nmos ( level=54                         lmin=1.8e-006                   lmax=9e-006 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.14344396 k2=0.013628333                minv=-0.4761                    cit=0.0001 voff=-0.097953042               eta0=0.042028419                etab=-0.028573274 u0=0.041150369                ua=-2.4698317e-011            ub=2.811627e-018 uc=1.8244874e-011             vsat=80000                      a0=8.034451 ags=0.93288333                 keta=-0.018167808               pclm=0.76297619 pdiblc2=0.0022540278               tvoff=0.00381828                 ltvoff=2.11358e-009 wtvoff=6.12986e-011               ptvoff=-5.80102e-016              kt1=-0.13386761 kt2=-0.021283821               ute=-1.7207464                 ua1=1.6314709e-009 ub1=-3.8484589e-018            uc1=-3.3831269e-011            at=75529.928 lvth0=2.8005279e-008             lk2=-7.7657619e-009            lvoff=1.4628754e-008 leta0=2.2943588e-007             lu0=2.950666e-009              lua=8.6075381e-017 lub=-3.2357341e-025            luc=2.5957658e-017             la0=-6.7461174e-006 lags=1.1221526e-006             lketa=-6.1236268e-008            lpclm=2.1355845e-006 lpdiblc2=-7.4421885e-010            lkt1=-2.6613913e-008            lkt2=5.1923017e-008 lute=5.8210857e-008             lua1=-6.5154742e-016            lub1=-1.1943095e-025 luc1=-4.1030403e-017            lat=-0.0047746493              letab=3.7503793e-007 lvsat=0                          lcit=0                          wvth0=6.922125e-009 wk2=-4.7331e-009               wvoff=3.740145e-009              weta0=5.5192071e-009 wu0=3.4327821e-010             wua=2.2718832e-017             wub=-2.1220714e-025 wuc=1.1555874e-017             wa0=-1.4879404e-006            wags=-3.8949e-008 wketa=1.1448482e-008             wpdiblc2=-7.365e-010                wkt1=-2.5507982e-008 wkt2=6.2238466e-009             wute=-4.4544429e-008            wua1=-4.0173193e-016 wub1=6.5689832e-025             wuc1=-7.3328764e-018            wat=0.0003271575 pvth0=-1.3366818e-014            pk2=1.5725668e-014             pvoff=-4.7599849e-014 peta0=-4.9728056e-014            pu0=-9.31309e-016              pua=-2.7158228e-023 pub=1.0483779e-031             puc=1.5104731e-023             pa0=8.9531469e-013 pags=-1.3279453e-014            pketa=-3.5382753e-014            wpclm=3.8785714e-008 ppclm=-3.4945929e-013            ppdiblc2=5.9408079e-015             pkt1=4.2808763e-015 pkt2=-5.6076858e-014            pute=5.381673e-014              pua1=2.6873419e-022 pub1=-4.527245e-031             puc1=4.1617106e-023             pat=-2.9476891e-009 wetab=6.8392608e-009             petab=-9.1313886e-014            wvsat=0 pvsat=0                          wcit=0                          pcit=0 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.15 nmos ( level=54                         lmin=1.08e-006                  lmax=1.8e-006 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.14760873 k2=0.027789459                minv=-0.4761                    cit=-0.00082390476 voff=-0.12172654                eta0=0.27400817                 etab=0.40296346 u0=0.041542643                ua=4.3790476e-012             ub=2.8216607e-018 uc=9.2651253e-011             vsat=81297.619                  a0=3.6695778 ags=1.4468849                  keta=-0.064543651               pclm=3.9109127 pdiblc2=-0.004282121               tvoff=0.00521724                 ltvoff=-4.18537e-010 wtvoff=-2.07931e-010              ptvoff=-9.27968e-017              kt1=-0.14986905 kt2=0.007634878                ute=-1.7175875                 ua1=1.5074547e-009 ub1=-4.532023e-018             uc1=-8.1053115e-011            at=135534.13 lvth0=3.5543516e-008             lk2=-3.33974e-008              lvoff=5.7658785e-008 leta0=-1.9044748e-007            lu0=2.2406507e-009             lua=3.3445352e-017 lub=-3.4173446e-025            luc=-1.0871789e-016            la0=1.1543031e-006 lags=1.9180972e-007             lketa=2.2704008e-008             lpclm=-3.5621806e-006 lpdiblc2=1.1086211e-008             lkt1=2.3486905e-009             lkt2=-4.1982842e-010 lute=5.2493232e-008             lua1=-4.2707805e-016            lub1=1.1178201e-024 luc1=4.4441138e-017             lat=-0.11338225                letab=-4.0604357e-007 lvsat=-0.0023486905              lcit=1.6722676e-009             wvth0=1.1098929e-008 wk2=-5.3451161e-009            wvoff=-1.4105571e-009            weta0=-7.2709929e-008 wu0=-2.2731429e-010            wua=2.7670629e-017             wub=-2.1104357e-025 wuc=-4.0877729e-018            wa0=-9.7881e-007               wags=2.8071429e-007 wketa=1.1169643e-008             wpdiblc2=8.9971907e-009             wkt1=-2.1214286e-009 wkt2=-2.5008348e-008            wute=4.79025e-008               wua1=-1.7616975e-016 wub1=3.0890786e-025             wuc1=1.5297964e-017             wat=-0.0049381071 pvth0=-2.0926832e-014            pk2=1.6833417e-014             pvoff=-3.8277078e-014 peta0=9.1866679e-014             pu0=1.0146343e-016             pua=-3.6120981e-023 pub=1.0273172e-031             puc=4.3419731e-023             pa0=-2.6211386e-014 pags=-5.9187e-013               pketa=-3.4878054e-014            wpclm=-9.7178571e-007 ppclm=1.479675e-012              ppdiblc2=-1.1677172e-014            pkt1=-3.8048786e-014 pkt2=4.534147e-016              pute=-1.1351221e-013            pua1=-1.3953335e-022 pub1=1.7713824e-031             puc1=6.5528464e-025             pat=6.5824399e-009 wetab=-1.2525179e-007            petab=1.4777092e-013             wvsat=-0.0014014286 pvsat=2.5365857e-009             wcit=2.1138214e-010             pcit=-3.8260168e-016 lmin_flag=1                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.model nch_na18ud15_mac.16 nmos ( level=54                         lmin=7.2e-07                    lmax=1.08e-006 wmin=4.5e-07                    wmax=1.08e-006                  vth0=-0.095765079 k2=-0.03964004                minv=-1.1083901                 cit=-0.00065133809 voff=0.081284921                eta0=0.16330556                 etab=0.059083575 u0=0.043725167                ua=5.9813333e-011             ub=3.051877e-018 uc=-6.376962e-011             vsat=76018.921                  a0=10.247024 ags=2.3325794                  keta=0.017119048                pclm=-0.081349206 pdiblc2=0.016091623                tvoff=0.00485724                 ltvoff=-2.61444e-011 wtvoff=-2.37341e-009              ptvoff=2.26757e-015               kt1=-0.11411111 kt2=0.076537722                ute=-1.5808147                 ua1=1.8498085e-009 ub1=-4.9514365e-018            uc1=-1.5588913e-010            at=74673.516 lvth0=-2.0966063e-008            lk2=4.0100754e-008             lvoff=-1.6362371e-007 leta0=-6.9781627e-008            lu0=-1.3830024e-010            lua=-2.6978019e-017 lub=-5.926702e-025             luc=6.1780863e-017             la0=-6.0151131e-006 lags=-7.7359722e-007            lketa=-6.6308333e-008            lpclm=7.8938492e-007 lpdiblc2=-1.1121171e-008            lkt1=-3.662746e-008             lkt2=-7.5523929e-008 lute=-9.6589139e-008            lua1=-8.002437e-016             lub1=1.5749808e-024 luc1=1.2601239e-016             lat=-0.047044184               letab=-3.121449e-008 lvsat=0.0034050908               lminv=6.8919619e-007             lcit=1.4841699e-009 wvth0=-2.0770714e-008            wk2=2.5741243e-008             wminv=7.8214286e-008 wvoff=-9.4953214e-008            weta0=2.565e-008                 wu0=-1.9707e-009 wua=-3.21984e-017              wub=-4.0837714e-025            wuc=5.2895919e-017 wa0=-3.4587857e-006            wags=-4.8128571e-007            wketa=-5.3678571e-008 wpdiblc2=-5.5079529e-009            wkt1=-3.9375e-008               wkt2=-2.5487925e-008 wute=-1.1317714e-007            wua1=-8.6719971e-016            wub1=1.3749514e-024 wuc1=-8.46786e-019              wat=-0.0057194571              pvth0=1.3811079e-014 pk2=-1.7050714e-014            pminv=-8.5253571e-014            pvoff=6.3684418e-014 peta0=-1.5345643e-014            pu0=2.0017539e-015             pua=2.9136261e-023 pub=3.1782531e-031             puc=-1.8692494e-023            pa0=2.6769621e-012 pags=2.3871e-013                pketa=3.58065e-014               wpclm=1.1678571e-006 ppclm=-8.5253571e-013            ppdiblc2=4.1334342e-015             pkt1=2.5576071e-015 pkt2=9.7615339e-016             pute=6.20646e-014               pua1=6.1368931e-022 pub1=-9.8484926e-031            puc1=1.8253063e-023             pat=7.4341114e-009 wetab=2.8732629e-008             petab=-2.0072101e-014            wvsat=0.0032439857 pvsat=-2.5269159e-009            wcit=-7.4397857e-011            pcit=-7.1101479e-017 lmin_flag=0                          lmax_flag=1                          wmin_flag=0 wmax_flag=1 tmimodel=1 )
.param random_fn_c=agauss(0,1,1) random_fn_io=agauss(0,1,1) r1_c=agauss(0,1,1) r2_c=agauss(0,1,1) r3_c=agauss(0,1,1) r4_c=agauss(0,1,1) r5_c=agauss(0,1,1) par1=r1_c par2=r2_c par3=r3_c par4=r4_c par5=r5_c r6_c=agauss(0,1,1) r7_c=0             r8_c=0             r9_c=0             r10_c=0 par6=r6_c par7=r7_c par8=r8_c par9=r9_c par10=r10_c r11_c=agauss(0,1,1) r12_c=agauss(0,1,1) r13_c=agauss(0,1,1) r14_c=agauss(0,1,1) r15_c=agauss(0,1,1) par11=r11_c par12=r12_c par13=r13_c par14=r14_c par15=r15_c r16_c=agauss(0,1,1) r17_c=0             r18_c=0             r19_c=0             r20_c=0 par16=r16_c par17=r17_c par18=r18_c par19=r19_c par20=r20_c r21_c=agauss(0,1,1) r22_c=agauss(0,1,1) r23_c=agauss(0,1,1) r24_c=agauss(0,1,1) r25_c=agauss(0,1,1) par21=r21_c par22=r22_c par23=r23_c par24=r24_c par25=r25_c r26_c=agauss(0,1,1) r27_c=0             r28_c=0             r29_c=0             r30_c=0 par26=r26_c par27=r27_c par28=r28_c par29=r29_c par30=r30_c r31_c=agauss(0,1,1) r32_c=agauss(0,1,1) par31=r31_c par32=r32_c r1_io=agauss(0,1,1) r2_io=agauss(0,1,1) r3_io=0             r4_io=0             r5_io=0 par1_io=r1_io par2_io=r2_io par3_io=r3_io par4_io=r4_io par5_io=r5_io r6_io=0             r7_io=agauss(0,1,1) r8_io=agauss(0,1,1) r9_io=0             r10_io=0 par6_io=r6_io par7_io=r7_io par8_io=r8_io par9_io=r9_io par10_io=r10_io r11_io=0             r12_io=0             r13_io=agauss(0,1,1) r14_io=agauss(0,1,1) r15_io=0 par11_io=r11_io par12_io=r12_io par13_io=r13_io par14_io=r14_io par15_io=r15_io r16_io=0             r17_io=0             r18_io=0             r19_io=agauss(0,1,1) r20_io=agauss(0,1,1) par16_io=r16_io par17_io=r17_io par18_io=r18_io par19_io=r19_io par20_io=r20_io plo_tox=agauss(0,1,1) plo_dxl=agauss(0,1,1) plo_dxw=agauss(0,1,1) parl1=agauss(0,1,1) parl2=agauss(0,1,1) parl3=agauss(0,1,1) parl4=agauss(0,1,1) parl5=agauss(0,1,1) r1_cap=agauss(0,1,1) r2_cap=agauss(0,1,1) par1_cap=r1_cap par2_cap=r2_cap w1_c='2.3875*0.35355' w2_c='0.70711*-0.35355' w3_c='0.54772*-0.0052117' w4_c='0.54772*-0.40307' w5_c='0.54772*-0.64548' w6_c='0.54772*-0.049915' w7_c='0.54772*-0.11513' w8_c='0.54772*-0.39385' w9_c=0 w10_c=0 w11_c='2.3875*0.35355' w12_c='0.70711*0.35355' w13_c='0.54772*0.32451' w14_c='0.54772*-0.16328' w15_c='0.54772*0.12195' w16_c='0.54772*0.66871' w17_c='0.54772*0.32929' w18_c='0.54772*-0.21807' w19_c=0 w20_c=0 w21_c='2.3875*0.35355' w22_c='0.70711*-0.35355' w23_c='0.54772*0.0088697' w24_c='0.54772*-0.21218' w25_c='0.54772*0.7283' w26_c='0.54772*-0.28609' w27_c='0.54772*-0.0042275' w28_c='0.54772*-0.30433' w29_c=0 w30_c=0 w31_c='2.3875*0.35355' w32_c='0.70711*0.35355' w33_c='0.54772*0.31715' w34_c='0.54772*0.2225' w35_c='0.54772*-0.17742' w36_c='0.54772*-0.6346' w37_c='0.54772*0.40656' w38_c='0.54772*0.020451' w39_c=0 w40_c=0 w41_c='2.3875*0.35355' w42_c='0.70711*-0.35355' w43_c='0.54772*0.0021707' w44_c='0.54772*0.81882' w45_c='0.54772*-0.058492' w46_c='0.54772*0.23016' w47_c='0.54772*-0.11085' w48_c='0.54772*-0.10416' w49_c=0 w50_c=0 w51_c='2.3875*0.35355' w52_c='0.70711*0.35355' w53_c='0.54772*0.22143' w54_c='0.54772*-0.066279' w55_c='0.54772*0.050463' w56_c='0.54772*-0.03945' w57_c='0.54772*-0.80208' w58_c='0.54772*0.22166' w59_c=0 w60_c=0 w61_c='2.3875*0.35355' w62_c='0.70711*-0.35355' w63_c='0.54772*-0.0058287' w64_c='0.54772*-0.20357' w65_c='0.54772*-0.024322' w66_c='0.54772*0.10585' w67_c='0.54772*0.2302' w68_c='0.54772*0.80233' w69_c=0 w70_c=0 w71_c='2.3875*0.35355' w72_c='0.70711*0.35355' w73_c='0.54772*-0.86309' w74_c='0.54772*0.007054' w75_c='0.54772*0.0050038' w76_c='0.54772*0.0053387' w77_c='0.54772*0.066237' w78_c='0.54772*-0.024037' w79_c=0 w80_c=0 w81_c=0 w82_c=0 w83_c=0 w84_c=0 w85_c=0 w86_c=0 w87_c=0 w88_c=0 w89_c=0 w90_c=0 w91_c=0 w92_c=0 w93_c=0 w94_c=0 w95_c=0 w96_c=0 w97_c=0 w98_c=0 w99_c=0 w100_c=0 w1_io='2.0857*0.40825' w2_io='0.67082*-0.40825' w3_io='0.54772*0.26807' w4_io='0.54772*-0.6902' w5_io='0.54772*-0.32981' w6_io='0.54772*0.098267' w7_io='2.0857*0.40825' w8_io='0.67082*0.40825' w9_io='0.54772*-0.10446' w10_io='0.54772*0.14211' w11_io='0.54772*-0.14894' w12_io='0.54772*0.78318' w13_io='2.0857*0.40825' w14_io='0.67082*-0.40825' w15_io='0.54772*0.51125' w16_io='0.54772*0.62722' w17_io='0.54772*0.10605' w18_io='0.54772*-0.025445' w19_io='2.0857*0.40825' w20_io='0.67082*0.40825' w21_io='0.54772*-0.094515' w22_io='0.54772*0.148' w23_io='0.54772*-0.55665' w24_io='0.54772*-0.57094' w25_io='2.0857*0.40825' w26_io='0.67082*-0.40825' w27_io='0.54772*-0.77931' w28_io='0.54772*0.062984' w29_io='0.54772*0.22376' w30_io='0.54772*-0.072822' w31_io='2.0857*0.40825' w32_io='0.67082*0.40825' w33_io='0.54772*0.19898' w34_io='0.54772*-0.2901' w35_io='0.54772*0.7056' w36_io='0.54772*-0.21225' p1_c1n='w1_c*par1+w2_c*par2+w3_c*par3+w4_c*par4+w5_c*par5+w6_c*par6+w7_c*par7+w8_c*par8+w9_c*par9+w10_c*par10' p1_c1p='w11_c*par1+w12_c*par2+w13_c*par3+w14_c*par4+w15_c*par5+w16_c*par6+w17_c*par7+w18_c*par8+w19_c*par9+w20_c*par10' p1_c2n='w21_c*par1+w22_c*par2+w23_c*par3+w24_c*par4+w25_c*par5+w26_c*par6+w27_c*par7+w28_c*par8+w29_c*par9+w30_c*par10' p1_c2p='w31_c*par1+w32_c*par2+w33_c*par3+w34_c*par4+w35_c*par5+w36_c*par6+w37_c*par7+w38_c*par8+w39_c*par9+w40_c*par10' p1_c3n='w41_c*par1+w42_c*par2+w43_c*par3+w44_c*par4+w45_c*par5+w46_c*par6+w47_c*par7+w48_c*par8+w49_c*par9+w50_c*par10' p1_c3p='w51_c*par1+w52_c*par2+w53_c*par3+w54_c*par4+w55_c*par5+w56_c*par6+w57_c*par7+w58_c*par8+w59_c*par9+w60_c*par10' p1_c4n='w61_c*par1+w62_c*par2+w63_c*par3+w64_c*par4+w65_c*par5+w66_c*par6+w67_c*par7+w68_c*par8+w69_c*par9+w70_c*par10' p1_c4p='w71_c*par1+w72_c*par2+w73_c*par3+w74_c*par4+w75_c*par5+w76_c*par6+w77_c*par7+w78_c*par8+w79_c*par9+w80_c*par10' p1_c5n='w81_c*par1+w82_c*par2+w83_c*par3+w84_c*par4+w85_c*par5+w86_c*par6+w87_c*par7+w88_c*par8+w89_c*par9+w90_c*par10' p1_c5p='w91_c*par1+w92_c*par2+w93_c*par3+w94_c*par4+w95_c*par5+w96_c*par6+w97_c*par7+w98_c*par8+w99_c*par9+w100_c*par10' p2_c1n='w1_c*par11+w2_c*par12+w3_c*par13+w4_c*par14+w5_c*par15+w6_c*par16+w7_c*par17+w8_c*par18+w9_c*par19+w10_c*par20' p2_c1p='w11_c*par11+w12_c*par12+w13_c*par13+w14_c*par14+w15_c*par15+w16_c*par16+w17_c*par17+w18_c*par18+w19_c*par19+w20_c*par20' p2_c2n='w21_c*par11+w22_c*par12+w23_c*par13+w24_c*par14+w25_c*par15+w26_c*par16+w27_c*par17+w28_c*par18+w29_c*par19+w30_c*par20' p2_c2p='w31_c*par11+w32_c*par12+w33_c*par13+w34_c*par14+w35_c*par15+w36_c*par16+w37_c*par17+w38_c*par18+w39_c*par19+w40_c*par20' p2_c3n='w41_c*par11+w42_c*par12+w43_c*par13+w44_c*par14+w45_c*par15+w46_c*par16+w47_c*par17+w48_c*par18+w49_c*par19+w50_c*par20' p2_c3p='w51_c*par11+w52_c*par12+w53_c*par13+w54_c*par14+w55_c*par15+w56_c*par16+w57_c*par17+w58_c*par18+w59_c*par19+w60_c*par20' p2_c4n='w61_c*par11+w62_c*par12+w63_c*par13+w64_c*par14+w65_c*par15+w66_c*par16+w67_c*par17+w68_c*par18+w69_c*par19+w70_c*par20' p2_c4p='w71_c*par11+w72_c*par12+w73_c*par13+w74_c*par14+w75_c*par15+w76_c*par16+w77_c*par17+w78_c*par18+w79_c*par19+w80_c*par20' p2_c5n='w81_c*par11+w82_c*par12+w83_c*par13+w84_c*par14+w85_c*par15+w86_c*par16+w87_c*par17+w88_c*par18+w89_c*par19+w90_c*par20' p2_c5p='w91_c*par11+w92_c*par12+w93_c*par13+w94_c*par14+w95_c*par15+w96_c*par16+w97_c*par17+w98_c*par18+w99_c*par19+w100_c*par20' p3_c1n='w1_c*par21+w2_c*par22+w3_c*par23+w4_c*par24+w5_c*par25+w6_c*par26+w7_c*par27+w8_c*par28+w9_c*par29+w10_c*par30' p3_c1p='w11_c*par21+w12_c*par22+w13_c*par23+w14_c*par24+w15_c*par25+w16_c*par26+w17_c*par27+w18_c*par28+w19_c*par29+w20_c*par30' p3_c2n='w21_c*par21+w22_c*par22+w23_c*par23+w24_c*par24+w25_c*par25+w26_c*par26+w27_c*par27+w28_c*par28+w29_c*par29+w30_c*par30' p3_c2p='w31_c*par21+w32_c*par22+w33_c*par23+w34_c*par24+w35_c*par25+w36_c*par26+w37_c*par27+w38_c*par28+w39_c*par29+w40_c*par30' p3_c3n='w41_c*par21+w42_c*par22+w43_c*par23+w44_c*par24+w45_c*par25+w46_c*par26+w47_c*par27+w48_c*par28+w49_c*par29+w50_c*par30' p3_c3p='w51_c*par21+w52_c*par22+w53_c*par23+w54_c*par24+w55_c*par25+w56_c*par26+w57_c*par27+w58_c*par28+w59_c*par29+w60_c*par30' p3_c4n='w61_c*par21+w62_c*par22+w63_c*par23+w64_c*par24+w65_c*par25+w66_c*par26+w67_c*par27+w68_c*par28+w69_c*par29+w70_c*par30' p3_c4p='w71_c*par21+w72_c*par22+w73_c*par23+w74_c*par24+w75_c*par25+w76_c*par26+w77_c*par27+w78_c*par28+w79_c*par29+w80_c*par30' p3_c5n='w81_c*par21+w82_c*par22+w83_c*par23+w84_c*par24+w85_c*par25+w86_c*par26+w87_c*par27+w88_c*par28+w89_c*par29+w90_c*par30' p3_c5p='w91_c*par21+w92_c*par22+w93_c*par23+w94_c*par24+w95_c*par25+w96_c*par26+w97_c*par27+w98_c*par28+w99_c*par29+w100_c*par30' p4_c1n='par31' p4_c1p='par31' p4_c2n='par31' p4_c2p='par31' p4_c3n='par31' p4_c3p='par31' p4_c4n='par31' p4_c4p='par31' p4_c5n='par31' p4_c5p='par31' p5_c1n='par32' p5_c1p='par32' p5_c2n='par32' p5_c2p='par32' p5_c3n='par32' p5_c3p='par32' p5_c4n='par32' p5_c4p='par32' p5_c5n='par32' p5_c5p='par32' p1_io1n='w1_io*par1_io+w2_io*par2_io+w3_io*par3_io+w4_io*par4_io+w5_io*par5_io+w6_io*par6_io' p1_io1p='w7_io*par1_io+w8_io*par2_io+w9_io*par3_io+w10_io*par4_io+w11_io*par5_io+w12_io*par6_io' p1_io2n='w13_io*par1_io+w14_io*par2_io+w15_io*par3_io+w16_io*par4_io+w17_io*par5_io+w18_io*par6_io' p1_io2p='w19_io*par1_io+w20_io*par2_io+w21_io*par3_io+w22_io*par4_io+w23_io*par5_io+w24_io*par6_io' p1_io3n='w25_io*par1_io+w26_io*par2_io+w27_io*par3_io+w28_io*par4_io+w29_io*par5_io+w30_io*par6_io' p1_io3p='w31_io*par1_io+w32_io*par2_io+w33_io*par3_io+w34_io*par4_io+w35_io*par5_io+w36_io*par6_io' p2_io1n='w1_io*par7_io+w2_io*par8_io+w3_io*par9_io+w4_io*par10_io+w5_io*par11_io+w6_io*par12_io' p2_io1p='w7_io*par7_io+w8_io*par8_io+w9_io*par9_io+w10_io*par10_io+w11_io*par11_io+w12_io*par12_io' p2_io2n='w13_io*par7_io+w14_io*par8_io+w15_io*par9_io+w16_io*par10_io+w17_io*par11_io+w18_io*par12_io' p2_io2p='w19_io*par7_io+w20_io*par8_io+w21_io*par9_io+w22_io*par10_io+w23_io*par11_io+w24_io*par12_io' p2_io3n='w25_io*par7_io+w26_io*par8_io+w27_io*par9_io+w28_io*par10_io+w29_io*par11_io+w30_io*par12_io' p2_io3p='w31_io*par7_io+w32_io*par8_io+w33_io*par9_io+w34_io*par10_io+w35_io*par11_io+w36_io*par12_io' p3_io1n='w1_io*par13_io+w2_io*par14_io+w3_io*par15_io+w4_io*par16_io+w5_io*par17_io+w6_io*par18_io' p3_io1p='w7_io*par13_io+w8_io*par14_io+w9_io*par15_io+w10_io*par16_io+w11_io*par17_io+w12_io*par18_io' p3_io2n='w13_io*par13_io+w14_io*par14_io+w15_io*par15_io+w16_io*par16_io+w17_io*par17_io+w18_io*par18_io' p3_io2p='w19_io*par13_io+w20_io*par14_io+w21_io*par15_io+w22_io*par16_io+w23_io*par17_io+w24_io*par18_io' p3_io3n='w25_io*par13_io+w26_io*par14_io+w27_io*par15_io+w28_io*par16_io+w29_io*par17_io+w30_io*par18_io' p3_io3p='w31_io*par13_io+w32_io*par14_io+w33_io*par15_io+w34_io*par16_io+w35_io*par17_io+w36_io*par18_io' p4_io1n='par19_io' p4_io1p='par19_io' p4_io2n='par19_io' p4_io2p='par19_io' p4_io3n='par19_io' p4_io3p='par19_io' p5_io1n='par20_io' p5_io1p='par20_io' p5_io2n='par20_io' p5_io2p='par20_io' p5_io3n='par20_io' p5_io3p='par20_io' par1fn_mc_c='random_fn_c' par1fn_mc_io='random_fn_io'
.option geoshrink=0.9
.param mismatchflag_bip=1
.param par_bjtp1=agauss(0,1,1) par_bjtp2=agauss(0,1,1) bfa=1        isa=1        nfa=1        rba=1        rea=1 rca=1        rbma=1        cjea=1        cjca=1
.model pnp10 pnp (                                             level=1 is='5.62e-018*isa'      bf='0.742*bfa'          nf='1.002*nfa' vaf=500                  ikf=0.01                 ise='1.27e-015*isa' ne=1.55                 br=0.00744              nr=0.99 var=41.65                ikr=0.00161              isc='5.62e-018*isa' nc=1.0618               rb='61.6*rba'           irb=0.00681 rbm='3*rbma'             re='13.27*rea'          rc='38*rca' nkf=0.22                 subs=1                    tref=25 xtb=0                    xti=3.41                 eg=1.1646 tlev=1                    tlevc=1                    tbf1=0.0036598 tbf2=-4.0899e-006         tbr1=0.0005837            tbr2=9.9e-007 tikf1=-0.0061838           tne1=0.00045              tnf1=1.8911e-005 tnf2=-8.64e-008           tnr1=-0.00014233          trb1=0.0034068 trc1=0.00025              tre1=0.00027242           tvar1=1e-011 cje='1.494e-13*cjea'     vje=0.789                mje=0.432 cjc='3.249e-14*cjca'     vjc=0.51                 mjc=0.292 fc=0                    ctc=0.00128              cte=0.00076 tvjc=0.00186              tvje=0.00105              )
.model pnp5 pnp (                                              level=1 is='1.5e-018*isa'       bf='0.865*bfa'          nf='1.002*nfa' vaf=500                  ikf=0.0038               ise='6e-016*isa' ne=1.58                 br=0.00395              nr=0.972 var=41.65                ikr=0.0019               isc='1.5e-018*isa' nc=1.1475               rb='99.2*rba'           irb=0.0065 rbm='0.1*rbma'           re='11.38*rea'          rc='17*rca' nkf=0.22                 subs=1                    tref=25 xtb=0                    xti=3.57                 eg=1.1583 tlev=1                    tlevc=1                    tbf1=0.003832 tbf2=-3.9029e-006         tbr1=0.0011844            tikf1=-0.00645 tnc1=0.000115             tne1=0.0005               tnf1=1.1561e-005 tnf2=-1.8e-007            tnr1=-1e-005              trb1=0.0042452 trc1=0.001971             tre1=0.00022              cje='3.836e-14*cjea' vje=0.789                mje=0.432                cjc='1.414e-14*cjca' vjc=0.51                 mjc=0.292                fc=0 ctc=0.00128              cte=0.00076              tvjc=0.00186 tvje=0.00105              )
.model pnp2 pnp (                                              level=1 is='2.85e-019*isa'      bf='1.362*bfa'          nf='1.0025*nfa' vaf=800                  ikf=0.0007               ise='1.85e-016*isa' ne=1.6                  br=0.00167              nr=0.968 var=35.1                 ikr=0.0008               isc='2.85e-019*isa' nc=1.19                 rb='210*rba'            irb=0.0013 rbm='0.1*rbma'           re='24*rea'             rc='39.175*rca' nkf=0.23                 subs=1                    tref=25 xtb=0                    xti=3                    eg=1.1814 tlev=1                    tlevc=1                    tbf1=0.0039168 tbf2=-3.09e-006           tbr1=0.0016852            tikf1=-0.006 tikr1=-6.042e-012          tnc1=5.17e-005            tne1=0.000455 tnf1=5.6e-005             tnf2=-2.664e-007          tnr1=-0.00024 trb1=0.0026356            trc1=0.00024              tre1=0.00021149 cje='6.625e-15*cjea'     vje=0.789                mje=0.432 cjc='6.270e-15*cjca'     vjc=0.51                 mjc=0.292 fc=0                    ctc=0.00128              cte=0.00076 tvjc=0.00186              tvje=0.00105              )
.subckt pnp10_mis c b e mismatchflag='mismatchflag_bip' multi='1'
.param ismis10='1+0.575e-2*(1/sqrt(multi*10e-6*10e-6*1e12*0.81))*par_bjtp1*mismatchflag' bfmis10='1+0.702e-2*(1/sqrt(multi*10e-6*10e-6*1e12*0.81))*par_bjtp2*mismatchflag'
qin c b e pnp10 m=multi
.model pnp10 pnp (                                             level=1 is='5.62e-018*isa*ismis10'      bf='0.742*bfa*bfmis10'          nf='1.002*nfa' vaf=500                  ikf=0.01                 ise='1.27e-015*isa/bfmis10' ne=1.55                 br=0.00744              nr=0.99 var=41.65                ikr=0.00161              isc='5.62e-018*isa' nc=1.0618               rb='61.6*rba'           irb=0.00681 rbm='3*rbma'             re='13.27*rea'          rc='38*rca' nkf=0.22                 subs=1                    tref=25 xtb=0                    xti=3.41                 eg=1.1646 tlev=1                    tlevc=1                    tbf1=0.0036598 tbf2=-4.0899e-006         tbr1=0.0005837            tbr2=9.9e-007 tikf1=-0.0061838           tne1=0.00045              tnf1=1.8911e-005 tnf2=-8.64e-008           tnr1=-0.00014233          trb1=0.0034068 trc1=0.00025              tre1=0.00027242           tvar1=1e-011 cje='1.494e-13*cjea'     vje=0.789                mje=0.432 cjc='3.249e-14*cjca'     vjc=0.51                 mjc=0.292 fc=0                    ctc=0.00128              cte=0.00076 tvjc=0.00186              tvje=0.00105              )
.ends pnp10_mis
.subckt pnp5_mis c b e mismatchflag='mismatchflag_bip' multi='1'
.param ismis5='1+0.575e-2*(1/sqrt(multi*5e-6*5e-6*1e12*0.81))*par_bjtp1*mismatchflag' bfmis5='1+0.702e-2*(1/sqrt(multi*5e-6*5e-6*1e12*0.81))*par_bjtp2*mismatchflag'
qin c b e pnp5 m=multi
.model pnp5 pnp (                                              level=1 is='1.5e-018*isa*ismis5'       bf='0.865*bfa*bfmis5'          nf='1.002*nfa' vaf=500                  ikf=0.0038               ise='6e-016*isa/bfmis5' ne=1.58                 br=0.00395              nr=0.972 var=41.65                ikr=0.0019               isc='1.5e-018*isa' nc=1.1475               rb='99.2*rba'           irb=0.0065 rbm='0.1*rbma'           re='11.38*rea'          rc='17*rca' nkf=0.22                 subs=1                    tref=25 xtb=0                    xti=3.57                 eg=1.1583 tlev=1                    tlevc=1                    tbf1=0.003832 tbf2=-3.9029e-006         tbr1=0.0011844            tikf1=-0.00645 tnc1=0.000115             tne1=0.0005               tnf1=1.1561e-005 tnf2=-1.8e-007            tnr1=-1e-005              trb1=0.0042452 trc1=0.001971             tre1=0.00022              cje='3.836e-14*cjea' vje=0.789                mje=0.432                cjc='1.414e-14*cjca' vjc=0.51                 mjc=0.292                fc=0 ctc=0.00128              cte=0.00076              tvjc=0.00186 tvje=0.00105              )
.ends pnp5_mis
.subckt pnp2_mis c b e mismatchflag='mismatchflag_bip' multi='1'
.param ismis2='1+0.575e-2*(1/sqrt(multi*2e-6*2e-6*1e12*0.81))*par_bjtp1*mismatchflag' bfmis2='1+0.702e-2*(1/sqrt(multi*2e-6*2e-6*1e12*0.81))*par_bjtp2*mismatchflag'
qin c b e pnp2 m=multi
.model pnp2 pnp (                                              level=1 is='2.85e-019*isa*ismis2'      bf='1.362*bfa*bfmis2'          nf='1.0025*nfa' vaf=800                  ikf=0.0007               ise='1.85e-016*isa/bfmis2' ne=1.6                  br=0.00167              nr=0.968 var=35.1                 ikr=0.0008               isc='2.85e-019*isa' nc=1.19                 rb='210*rba'            irb=0.0013 rbm='0.1*rbma'           re='24*rea'             rc='39.175*rca' nkf=0.23                 subs=1                    tref=25 xtb=0                    xti=3                    eg=1.1814 tlev=1                    tlevc=1                    tbf1=0.0039168 tbf2=-3.09e-006           tbr1=0.0016852            tikf1=-0.006 tikr1=-6.042e-012          tnc1=5.17e-005            tne1=0.000455 tnf1=5.6e-005             tnf2=-2.664e-007          tnr1=-0.00024 trb1=0.0026356            trc1=0.00024              tre1=0.00021149 cje='6.625e-15*cjea'     vje=0.789                mje=0.432 cjc='6.270e-15*cjca'     vjc=0.51                 mjc=0.292 fc=0                    ctc=0.00128              cte=0.00076 tvjc=0.00186              tvje=0.00105              )
.ends pnp2_mis
.param mismatchflag_bip_npn=1
.param par_bjtn1=agauss(0,1,1) par_bjtn2=agauss(0,1,1) bfb=1        isb=1        nfb=1        rbb=1        reb=1 rcb=1        rbmb=1        cjeb=1        cjcb=1
.model npn10 npn (                                             level=1 is='9.75e-018*isb'      bf='5.69*bfb'           nf='0.9998*nfb' vaf=100                  ikf=0.02                 ise='1.0924e-016*isb' ne=1.4212               br=0.679                nr=0.995 var=39.602               ikr=0.0167               isc='9.75e-018*isb' nc=1.0753               rb='198.55*rbb'         irb=0.00056332 rbm='0.1*rbmb'           re='13.119*reb'         rc='12.358*rcb' nkf=0.2                  subs=1                    tref=25 xtb=0                    xti=3.604                eg=1.1625 tlev=1                    tlevc=1                    tbf1=0.003675 tbf2=-1.775e-006          tbr1=0.00078867           tbr2=-3e-006 tikf1=-0.00645             tikr1=1.71e-011            tne1=0.000472 tnf1=1.0739e-005          tnf2=-1e-007              tnr1=1e-005 trb1=0.00134              trc1=0.0018358            tre1=0.00027242 cje='1.195e-13*cjeb'     vje=0.672                mje=0.321 cjc='7.8051e-14*cjcb'    vjc=0.701                mjc=0.338 fc=0                    ctc=0.00104              cte=0.00072 tvjc=0.0015               tvje=0.00114              )
.model npn5 npn (                                              level=1 is='2.605e-018*isb'     bf='6.1*bfb'            nf='0.9998*nfb' vaf=96.792               ikf=0.02                 ise='4.472e-017*isb' ne=1.4082               br=0.3848               nr=0.995 var=35.497               ikr=0.02                 isc='2.605e-018*isb' nc=1.1                  rb='420.8*rbb'          irb=0.0001509 rbm='0.1*rbmb'           re='29.906*reb'         rc='6.4768*rcb' nkf=0.38                 subs=1                    tref=25 xtb=0                    xti=3.54                 eg=1.164 tlev=1                    tlevc=1                    tbf1=0.0035859 tbf2=-2.1795e-006         tbr1=0.0006563            tbr2=-3e-006 tikf1=-0.0057517           tikr1=1.71e-011            tne1=0.00026973 tnf1=1e-005               tnf2=-1.552e-007          tnr1=1.2107e-005 trb1=0.0014               trc1=0.0055               tre1=0.00027242 cje='3.084e-14*cjeb'     vje=0.672                mje=0.321 cjc='2.8259e-14*cjcb'    vjc=0.701                mjc=0.338 fc=0                    ctc=0.00104              cte=0.00072 tvjc=0.0015               tvje=0.00114              )
.model npn2 npn (                                              level=1 is='4.972e-019*isb'     bf='7.1*bfb'            nf='1.001*nfb' vaf=92.856               ikf=0.0012379            ise='1.003e-017*isb' ne=1.36                 br=0.1645               nr=0.992 var=32.85                ikr=0.0016922            isc='4.972e-019*isb' nc=1.0251               rb='465.26*rbb'         irb=0.0001913 rbm='0.1*rbmb'           re='26.148*reb'         rc='17.26*rcb' nkf=0.22                 subs=1                    tref=25 xtb=0                    xti=3                    eg=1.1775 tlev=1                    tlevc=1                    tbf1=0.00333 tbf2=-6e-007              tbr1=0.00054789           tbr2=-2.3504e-006 tikf1=-0.0049              tikr1=1.71e-011            tne1=0.0004 tnf1=1.54e-005            tnf2=-3e-007              tnr1=-4e-005 trb1=0.001715             trc1=0.0018358            tre1=0.00027242 cje='5.396e-15*cjeb'     vje=0.672                mje=0.321 cjc='1.0108e-14*cjcb'    vjc=0.701                mjc=0.338 fc=0                    ctc=0.00104              cte=0.00072 tvjc=0.0015               tvje=0.00114              )
.subckt npn10_mis c b e mismatchflag='mismatchflag_bip_npn' multi='1'
.param ismis10='1+0.174e-2*(1/sqrt(multi*10e-6*10e-6*1e12*0.81))*par_bjtn1*mismatchflag' bfmis10='1+1.485e-2*(1/sqrt(multi*10e-6*10e-6*1e12*0.81))*par_bjtn2*mismatchflag'
qin c b e npn10 m=multi
.model npn10 npn (                                             level=1 is='9.75e-018*isb*ismis10'      bf='5.69*bfb*bfmis10'           nf='0.9998*nfb' vaf=100                  ikf=0.02                 ise='1.0924e-016*isb/bfmis10' ne=1.4212               br=0.679                nr=0.995 var=39.602               ikr=0.0167               isc='9.75e-018*isb' nc=1.0753               rb='198.55*rbb'         irb=0.00056332 rbm='0.1*rbmb'           re='13.119*reb'         rc='12.358*rcb' nkf=0.2                  subs=1                    tref=25 xtb=0                    xti=3.604                eg=1.1625 tlev=1                    tlevc=1                    tbf1=0.003675 tbf2=-1.775e-006          tbr1=0.00078867           tbr2=-3e-006 tikf1=-0.00645             tikr1=1.71e-011            tne1=0.000472 tnf1=1.0739e-005          tnf2=-1e-007              tnr1=1e-005 trb1=0.00134              trc1=0.0018358            tre1=0.00027242 cje='1.195e-13*cjeb'     vje=0.672                mje=0.321 cjc='7.8051e-14*cjcb'     vjc=0.701                mjc=0.338 fc=0                    ctc=0.00104              cte=0.00072 tvjc=0.0015               tvje=0.00114              )
.ends npn10_mis
.subckt npn5_mis c b e mismatchflag='mismatchflag_bip_npn' multi='1'
.param ismis5='1+0.174e-2*(1/sqrt(multi*5e-6*5e-6*1e12*0.81))*par_bjtn1*mismatchflag' bfmis5='1+1.485e-2*(1/sqrt(multi*5e-6*5e-6*1e12*0.81))*par_bjtn2*mismatchflag'
qin c b e npn5 m=multi
.model npn5 npn (                                              level=1 is='2.605e-018*isb*ismis5'     bf='6.1*bfb*bfmis5'            nf='0.9998*nfb' vaf=96.792               ikf=0.02                 ise='4.472e-017*isb/bfmis5' ne=1.4082               br=0.3848               nr=0.995 var=35.497               ikr=0.02                 isc='2.605e-018*isb' nc=1.1                  rb='420.8*rbb'          irb=0.0001509 rbm='0.1*rbmb'           re='29.906*reb'         rc='6.4768*rcb' nkf=0.38                 subs=1                    tref=25 xtb=0                    xti=3.54                 eg=1.164 tlev=1                    tlevc=1                    tbf1=0.0035859 tbf2=-2.1795e-006         tbr1=0.0006563            tbr2=-3e-006 tikf1=-0.0057517           tikr1=1.71e-011            tne1=0.00026973 tnf1=1e-005               tnf2=-1.552e-007          tnr1=1.2107e-005 trb1=0.0014               trc1=0.0055               tre1=0.00027242 cje='3.084e-14*cjeb'     vje=0.672                mje=0.321 cjc='2.8259e-14*cjcb'     vjc=0.701                mjc=0.338 fc=0                    ctc=0.00104              cte=0.00072 tvjc=0.0015               tvje=0.00114              )
.ends npn5_mis
.subckt npn2_mis c b e mismatchflag='mismatchflag_bip_npn' multi='1'
.param ismis2='1+0.174e-2*(1/sqrt(multi*2e-6*2e-6*1e12*0.81))*par_bjtn1*mismatchflag' bfmis2='1+1.485e-2*(1/sqrt(multi*2e-6*2e-6*1e12*0.81))*par_bjtn2*mismatchflag'
qin c b e npn2 m=multi
.model npn2 npn (                                              level=1 is='4.972e-019*isb*ismis2'     bf='7.1*bfb*bfmis2'            nf='1.001*nfb' vaf=92.856               ikf=0.0012379            ise='1.003e-017*isb/bfmis2' ne=1.36                 br=0.1645               nr=0.992 var=32.85                ikr=0.0016922            isc='4.972e-019*isb' nc=1.0251               rb='465.26*rbb'         irb=0.0001913 rbm='0.1*rbmb'           re='26.148*reb'         rc='17.26*rcb' nkf=0.22                 subs=1                    tref=25 xtb=0                    xti=3                    eg=1.1775 tlev=1                    tlevc=1                    tbf1=0.00333 tbf2=-6e-007              tbr1=0.00054789           tbr2=-2.3504e-006 tikf1=-0.0049              tikr1=1.71e-011            tne1=0.0004 tnf1=1.54e-005            tnf2=-3e-007              tnr1=-4e-005 trb1=0.001715             trc1=0.0018358            tre1=0.00027242 cje='5.396e-15*cjeb'     vje=0.672                mje=0.321 cjc='1.0108e-14*cjcb'     vjc=0.701                mjc=0.338 fc=0                    ctc=0.00104              cte=0.00072 tvjc=0.0015               tvje=0.00114              )
.ends npn2_mis
.param is_d=1         x_jsw_d=0         n_d=1         rs_d=1 cj_d=1         cjsw_d=1
.model ndio d (                                             level=3 n='1.03*n_d'           is='4.32e-07*is_d'         jsw='1.17e-13*pwr(2,x_jsw_d)' bv=8.219999                    tcv=-5.51e-04                   rs='1.0e-10*rs_d' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.428e-03*cj_d'       pb=0.672                        mj=0.321 cta=0.00072                   tpb=0.00114                    cjsw='1.069e-10*cjsw_d' php=0.480                    mjsw=0.016                       ctp=0.00020 tphp=0.00244                 jtun='1.69e-05*is_d'         jtunsw='5.06e-11*pwr(2,x_jsw_d)' ntun=42.17                     keg=0.45                        xtitun=3 xti=3.00                        eg=1.08                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model pdio d (                                             level=3 n='1.02*n_d'           is='4.45e-07*is_d'         jsw='9.12e-14*pwr(2,x_jsw_d)' bv=7.43                    tcv=-3.06e-04                   rs='1.0e-10*rs_d' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.794e-03*cj_d'       pb=0.789                        mj=0.432 cta=0.00076                   tpb=0.00105                    cjsw='1.129e-10*cjsw_d' php=0.770                    mjsw=0.277                       ctp=0.00034 tphp=0.00097                 jtun='5.22e-05*is_d'         jtunsw='1.52e-10*pwr(2,x_jsw_d)' ntun=28.76                     keg=0.41                        xtitun=3 xti=3.00                        eg=1.10                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model nwdio d (                                             level=3 n='1.02*n_d'           is='2.57e-06*is_d'         jsw='3.63e-13*pwr(2,x_jsw_d)' bv=14.93                    tcv=-1.26e-03                   rs='1.0e-10*rs_d' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.611e-04*cj_d'       pb=0.510                        mj=0.292 cta=0.00128                  tpb=0.00186                    cjsw='3.637e-10*cjsw_d' php=0.780                    mjsw=0.358                       ctp=0.00102 tphp=0.00196                 jtun='3.43e-09*is_d'         jtunsw='1e-12*pwr(2,x_jsw_d)' ntun=58.02                     keg=0.41                        xtitun=3 xti=3.00                        eg=1.10                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.000484                   area=1.4241e-08                       )
.param is_d_12=1         x_jsw_d_12=0         n_d_12=1         rs_d_12=1 cj_d_12=1         cjsw_d_12=1
.model ndio_12 d (                                             level=3 n='1.02*n_d_12'           is='2.24e-07*is_d_12'         jsw='7.31e-14*pwr(2,x_jsw_d_12)' bv=8.22                    tcv=-5.01e-04                   rs='1.0e-10*rs_d_12' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.44e-03*cj_d_12'       pb=0.672                        mj=0.327 cta=0.0008                   tpb=0.0013                    cjsw='1.13e-10*cjsw_d_12' php=0.438                    mjsw=0.008                       ctp=0.00016 tphp=0.00218                 jtun='2.88e-05*is_d_12'         jtunsw='5.66e-11*pwr(2,x_jsw_d_12)' ntun=46.88                     keg=0.45                        xtitun=3 xti=3.00                        eg=1.15                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model pdio_12 d (                                             level=3 n='1.02*n_d_12'           is='4.90e-07*is_d_12'         jsw='1.01e-13*pwr(2,x_jsw_d_12)' bv=7.42                    tcv=-5.13e-04                   rs='1.0e-10*rs_d_12' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.878e-03*cj_d_12'       pb=0.816                        mj=0.449 cta=0.00075                   tpb=0.00100                    cjsw='1.13e-10*cjsw_d_12' php=0.742                    mjsw=0.253                       ctp=0.00041 tphp=0.00098                 jtun='2.25e-05*is_d_12'         jtunsw='8.98e-11*pwr(2,x_jsw_d_12)' ntun=26.31                     keg=0.44                        xtitun=3 xti=3.00                        eg=1.10                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_18=1         x_jsw_d_18=0         n_d_18=1         rs_d_18=1 cj_d_18=1         cjsw_d_18=1
.model ndio_18 d (                                             level=3 n='1.09*n_d_18'           is='2.69e-07*is_d_18'         jsw='7.06e-14*pwr(2,x_jsw_d_18)' bv=7.9                    tcv=0.00e+00                   rs='1.0e-10*rs_d_18' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.472e-03*cj_d_18'       pb=0.715                        mj=0.336 cta=0.00079                   tpb=0.00137                    cjsw='1.086e-10*cjsw_d_18' php=0.457                    mjsw=0.015                       ctp=0.00020 tphp=0.00230                 jtun='1.93e-03*is_d_18'         jtunsw='1.67e-10*pwr(2,x_jsw_d_18)' ntun=33.83                     keg=0.29                        xtitun=3 xti=3.00                        eg=1.27                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model pdio_18 d (                                             level=3 n='1.02*n_d_18'           is='2.81e-07*is_d_18'         jsw='4.79e-14*pwr(2,x_jsw_d_18)' bv=7.34                    tcv=-2.42e-04                   rs='1.0e-10*rs_d_18' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.836e-03*cj_d_18'       pb=0.830                        mj=0.451 cta=0.00085                   tpb=0.00129                    cjsw='1.454e-10*cjsw_d_18' php=0.924                    mjsw=0.560                       ctp=0.00066 tphp=0.00107                 jtun='3.53e-05*is_d_18'         jtunsw='3.35e-11*pwr(2,x_jsw_d_18)' ntun=28.61                     keg=0.41                        xtitun=3 xti=3.00                        eg=1.13                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_18ud15=1         x_jsw_d_18ud15=0         n_d_18ud15=1         rs_d_18ud15=1 cj_d_18ud15=1         cjsw_d_18ud15=1
.model ndio_18ud15 d (                                             level=3 n='1.09*n_d_18ud15'           is='2.69e-07*is_d_18ud15'         jsw='7.06e-14*pwr(2,x_jsw_d_18ud15)' bv=7.9                    tcv=0.00e+00                   rs='1.0e-10*rs_d_18ud15' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.472e-03*cj_d_18ud15'       pb=0.715                        mj=0.336 cta=0.00079                   tpb=0.00137                    cjsw='1.086e-10*cjsw_d_18ud15' php=0.457                    mjsw=0.015                       ctp=0.00020 tphp=0.00230                 jtun='1.93e-03*is_d_18ud15'         jtunsw='1.67e-10*pwr(2,x_jsw_d_18ud15)' ntun=33.83                     keg=0.29                        xtitun=3 xti=3.00                        eg=1.27                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model pdio_18ud15 d (                                             level=3 n='1.02*n_d_18ud15'           is='2.81e-07*is_d_18ud15'         jsw='4.79e-14*pwr(2,x_jsw_d_18ud15)' bv=7.34                    tcv=-2.42e-04                   rs='1.0e-10*rs_d_18ud15' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.836e-03*cj_d_18ud15'       pb=0.830                        mj=0.451 cta=0.00085                   tpb=0.00129                    cjsw='1.454e-10*cjsw_d_18ud15' php=0.924                    mjsw=0.560                       ctp=0.00066 tphp=0.00107                 jtun='3.53e-05*is_d_18ud15'         jtunsw='3.35e-11*pwr(2,x_jsw_d_18ud15)' ntun=28.61                     keg=0.41                        xtitun=3 xti=3.00                        eg=1.13                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_dnw=1         x_jsw_d_dnw=0         n_d_dnw=1         rs_d_dnw=1 cj_d_dnw=1         cjsw_d_dnw=1
.model dnwpsub d (                                             level=3 n='1.068*n_d_dnw'           is='3.35e-06*is_d_dnw'         jsw='7.46e-12*pwr(2,x_jsw_d_dnw)' bv=14.64                    tcv=-8.65e-04                   rs='1.0e-10*rs_d_dnw' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.223e-04*cj_d_dnw'       pb=0.5200                        mj=0.3 cta=0.00070                   tpb=0.00117                    cjsw='9.339e-10*cjsw_d_dnw' php=0.5480                    mjsw=0.2417                       ctp=0.00058 tphp=0.00127                 jtun='1.48e-06*is_d_dnw'         jtunsw='1.19e-10*pwr(2,x_jsw_d_dnw)' ntun=239.40                     keg=0.60                        xtitun=3 xti=3.00                        eg=1.17                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.000484                   area=1.4241e-08                       )
.model pwdnw d (                                             level=3 n='0.997*n_d_dnw'           is='8.67e-08*is_d_dnw'         jsw='5.38e-14*pwr(2,x_jsw_d_dnw)' bv=14.95                    tcv=-1.21e-03                   rs='1.0e-10*rs_d_dnw' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='6.031e-04*cj_d_dnw'       pb=0.7010                        mj=0.338 cta=0.00104                   tpb=0.0015                    cjsw='3.128e-10*cjsw_d_dnw' php=0.7150                    mjsw=0.3597                       ctp=0.00125 tphp=0.0022                 jtun='2.55e-08*is_d_dnw'         jtunsw='2.38e-12*pwr(2,x_jsw_d_dnw)' ntun=68.35                     keg=0.72                        xtitun=3 xti=3.00                        eg=1.20                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_esd=1.0     x_jsw_d_esd=0      n_d_esd=1.000 rs_d_esd=1.0     cj_d_esd=1.00     cjsw_d_esd=1.00
.model ndio_esd d (  is='1.51e-07*is_d_esd'    jsw='6.21e-13*pwr(2,x_jsw_d_esd)'  rs='1.0e-10*rs_d_esd'     n='1.005*n_d_esd'  cj='1.57e-03*cj_d_esd'    cjsw='1.71e-10*cjsw_d_esd'  bv=7.20e+00               area=1.4e-8          pj=4.8e-4  mj=0.29                   mjsw=0.06            pb=0.7  php=0.25                   trs=2.5e-3          tcv=-5.56e-04  cta=7.44e-04               ctp=3.00e-04        tpb=1.40e-03  tphp=8.00e-04               ik=1e20            ikr=1e10  ibv=0.03                   tref=25              fc=0  fcs=0                      tlev=1               tlevc=1  xti=3                      eg=1.17            level=3  )
.param is_d_hvt=1         x_jsw_d_hvt=0         n_d_hvt=1         rs_d_hvt=1 cj_d_hvt=1         cjsw_d_hvt=1
.model ndio_hvt d (                                             level=3 n='1.02*n_d_hvt'           is='2.20e-07*is_d_hvt'         jsw='6.35e-14*pwr(2,x_jsw_d_hvt)' bv=8.02                    tcv=-3.22e-04                   rs='1.0e-10*rs_d_hvt' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.686e-03*cj_d_hvt' cjsw='1.31e-10*cjsw_d_hvt' pb=0.748                        mj=0.406 cta=0.00075                   tpb=0.00103 php=0.616                    mjsw=0.110                       ctp=0.00016 tphp=0.00067                 jtun='3.97e-05*is_d_hvt'         jtunsw='4.66e-11*pwr(2,x_jsw_d_hvt)' ntun=35.02                     keg=0.44                        xtitun=3 xti=3.00                        eg=1.15                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model pdio_hvt d (                                             level=3 n='1.02*n_d_hvt'           is='8.95e-07*is_d_hvt'         jsw='2.11e-13*pwr(2,x_jsw_d_hvt)' bv=7.0                    tcv=0.00e+00                   rs='1.0e-10*rs_d_hvt' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='2.426e-03*cj_d_hvt' cjsw='1.242e-10*cjsw_d_hvt' pb=0.938                        mj=0.518 cta=0.00069                   tpb=0.00096 php=0.777                    mjsw=0.253                       ctp=0.00021 tphp=0.00061                 jtun='1.11e-04*is_d_hvt'         jtunsw='1.33e-10*pwr(2,x_jsw_d_hvt)' ntun=20.00                     keg=0.45                        xtitun=3 xti=3.00                        eg=1.05                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_lvt=1         x_jsw_d_lvt=0         n_d_lvt=1         rs_d_lvt=1 cj_d_lvt=1         cjsw_d_lvt=1
.model ndio_lvt d (                                             level=3 n='1.03*n_d_lvt'           is='3.11e-07*is_d_lvt'         jsw='9.46e-14*pwr(2,x_jsw_d_lvt)' bv=8.32                    tcv=-4.84e-04                   rs='1.0e-10*rs_d_lvt' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.39e-03*cj_d_lvt'       pb=0.67                        mj=0.313 cta=0.00073                   tpb=0.00113                    cjsw='1.05e-10*cjsw_d_lvt' php=0.472                    mjsw=0.011                       ctp=0.00016 tphp=0.00240                 jtun='5.73e-06*is_d_lvt'         jtunsw='2.21e-11*pwr(2,x_jsw_d_lvt)' ntun=37.72                     keg=0.48                        xtitun=3 xti=3.00                        eg=1.14                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.model pdio_lvt d (                                             level=3 n='1.02*n_d_lvt'           is='3.97e-07*is_d_lvt'         jsw='8.37e-14*pwr(2,x_jsw_d_lvt)' bv=7.58                    tcv=-3.41e-04                   rs='1.0e-10*rs_d_lvt' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.73e-03*cj_d_lvt'       pb=0.778                        mj=0.421 cta=0.00079                   tpb=0.00104                    cjsw='1.07e-10*cjsw_d_lvt' php=0.751                    mjsw=0.254                       ctp=0.00030 tphp=0.00089                 jtun='2.40e-05*is_d_lvt'         jtunsw='3.40e-11*pwr(2,x_jsw_d_lvt)' ntun=27.73                     keg=0.46                        xtitun=3 xti=3.00                        eg=1.11                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_na=1         x_jsw_d_na=0         n_d_na=1         rs_d_na=1 cj_d_na=1         cjsw_d_na=1
.model ndio_na d (                                             level=3 n='1.02*n_d_na'           is='2.76e-06*is_d_na'         jsw='2.63e-12*pwr(2,x_jsw_d_na)' bv=17.22                    tcv=-5.5e-04                   rs='1.0e-10*rs_d_na' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.59e-04*cj_d_na'       pb=0.530                        mj=0.336 cta=0.0022                   tpb=0.0023                    cjsw='1.99e-10*cjsw_d_na' php=0.4                    mjsw=0.039                       ctp=0.00044 tphp=0.0019                 jtun='4.93e-04*is_d_na'                    jtunsw='1.00e-14*pwr(2,x_jsw_d_na)' ntun=234.06                     keg=0.45                        xtitun=3 xti=3.00                        eg=1.09                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_na12=1         x_jsw_d_na12=0         n_d_na12=1         rs_d_na12=1 cj_d_na12=1         cjsw_d_na12=1
.model ndio_na12 d (                                             level=3 n='1.02*n_d_na12'           is='1.28e-06*is_d_na12'         jsw='1.24e-12*pwr(2,x_jsw_d_na12)' bv=16.56                    tcv=-7.5e-04                   rs='1.0e-10*rs_d_na12' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.576e-04*cj_d_na12'       pb=0.542                        mj=0.340 cta=0.0023                   tpb=0.0023                    cjsw='2.102e-10*cjsw_d_na12' php=0.463                    mjsw=0.045                       ctp=0.00025 tphp=0.0018                 jtun='1.16e-04*is_d_na12'         jtunsw='7.57e-10*pwr(2,x_jsw_d_na12)' ntun=800                     keg=0.52                        xtitun=3 xti=3.00                        eg=1.17                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_na18=1         x_jsw_d_na18=0         n_d_na18=1         rs_d_na18=1 cj_d_na18=1         cjsw_d_na18=1
.model ndio_na18 d (                                             level=3 n='1.02*n_d_na18'           is='1.60e-06*is_d_na18'         jsw='1.57e-12*pwr(2,x_jsw_d_na18)' bv=19.65                    tcv=-5.8e-04                   rs='1.0e-10*rs_d_na18' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.61e-04*cj_d_na18'       pb=0.512                        mj=0.292 cta=0.0012                   tpb=0.0014                    cjsw='2.08e-10*cjsw_d_na18' php=0.3                    mjsw=0.039                       ctp=0.00034 tphp=0.0013                 jtun='4.66e-05*is_d_na18'         jtunsw='3.35e-10*pwr(2,x_jsw_d_na18)' ntun=900                     keg=0.55                        xtitun=3 xti=3.00                        eg=1.15                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param is_d_na18ud15=1         x_jsw_d_na18ud15=0         n_d_na18ud15=1         rs_d_na18ud15=1 cj_d_na18ud15=1         cjsw_d_na18ud15=1
.model ndio_na18ud15 d (                                             level=3 n='1.02*n_d_na18ud15'           is='1.60e-06*is_d_na18ud15'         jsw='1.57e-12*pwr(2,x_jsw_d_na18ud15)' bv=19.65                    tcv=-5.8e-04                   rs='1.0e-10*rs_d_na18ud15' ikr=1e10                     ibv=0.03                        trs=2.5e-3 cj='1.61e-04*cj_d_na18ud15'       pb=0.512                        mj=0.292 cta=0.0012                   tpb=0.0014                    cjsw='2.08e-10*cjsw_d_na18ud15' php=0.3                    mjsw=0.039                       ctp=0.00034 tphp=0.0013                 jtun='4.66e-05*is_d_na18ud15'         jtunsw='3.35e-10*pwr(2,x_jsw_d_na18ud15)' ntun=900                     keg=0.55                        xtitun=3 xti=3.00                        eg=1.15                        fc=0 fcs=0                        ik=1e20                        tref=25 tlev=1                        tlevc=1 pj=0.00048                   area=1.4e-08                       )
.param mismatchflag_disres=1 scale_disres=0.9 rnoiseflag_disres=0
.param par_disres=agauss(0,1,1) r_rnodwo_m=1.0930e+002       rend_rnodwo_m=9.5824e-006         x_dxw_rnodwo_m=0            dxl_rnodwo_m=0 r_rpodwo_m=3.1373e+002       rend_rpodwo_m=6.0000e-006         x_dxw_rpodwo_m=0            dxl_rpodwo_m=0 r_rnpolywo_m=1.4970e+002   rend_rnpolywo_m=7.5700e-006     x_dxw_rnpolywo_m=0        dxl_rnpolywo_m=0 r_rppolywo_m=8.7600e+002   rend_rppolywo_m=6.2372e-006     x_dxw_rppolywo_m=0        dxl_rppolywo_m=0 r_rnodl_m=1.8000e+001        dxl_rnodl_m=0                     x_dxw_rnodl_m=0 r_rnods_m=1.8000e+001        dxl_rnods_m=0                     x_dxw_rnods_m=0 r_rpodl_m=1.6700e+001        dxl_rpodl_m=0                     x_dxw_rpodl_m=0 r_rpods_m=1.6700e+001        dxl_rpods_m=0                     x_dxw_rpods_m=0 r_rnpolyl_m=1.6420e+001    dxl_rnpolyl_m=0                 x_dxw_rnpolyl_m=0 r_rnpolys_m=1.6420e+001    dxl_rnpolys_m=0                 x_dxw_rnpolys_m=0 r_rppolyl_m=1.4400e+001    dxl_rppolyl_m=0                 x_dxw_rppolyl_m=0 r_rppolys_m=1.4400e+001    dxl_rppolys_m=0                 x_dxw_rppolys_m=0 r_rnwod_m=385                           rend_rnwod_m='170e-6' r_rnwsti_m=1169                        rend_rnwsti_m='2.7e-4' ca_pofox=1.079e-16                     cf_posfox=3.73e-17              cf_polfox=4.87e-17 ca_pofox_r=1.079e-16                    cf_polfox_r=4.87e-17
.subckt rnodwo_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00198323903818953*geo_fac*par_disres*mismatchflag'
.param rsh='r_rnodwo_m'     rendsh='2*rend_rnodwo_m*1e6'
.param dw_etch='0-9.25714285714286e-08*(pwr(0.5625,x_dxw_rnodwo_m)-1)'
.param dw_emp='1.5370e-009'     dw_empend='-5.2360e-008'
.param dl_etch='0+dxl_rnodwo_m'     dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'     dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=0.411133860400214
.param jc1_w=0.0577271204979308     jc1_n=-0.00313
.param jc1end_0=-1.13929     jc1end_w=40.82881
.param tc1_0=0.0014342814911298     tc1_w=-2.24331695355166e-07
.param tc2_0=7.54746914856436e-07     tc2_w=-2.0217e-09
.param tc1end_0=0.00135719397917256     tc1end_w=2.1275e-05
.param tc2end_0=3.37552662511097e-07     tc2end_w=-1.481e-08
.param jct_0=-0.00027337     jct_w=0.00019370448410292
.param jct_n=-3.8271e-06     jctend_0=-0.0487
.param jctend_w=0.0962829566646918     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 25)'
.param tc2='tc2_0 + tc2_w * min(wum, 25)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 25)'
.param tc2end='tc2end_0 + tc2end_w * min(wum, 25)'
.param jct='jct_0 + jct_w * min(wum, 25) + jct_n * min(nsqr, 150)'
.param jctend='jctend_0 + jctend_w * min(wum, 25)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 25) + jc1_n * min(nsqr, 150) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param jc1end='max(0, (jc1end_0 + jc1end_w * min(wum, 25) + jctend * delta_t))'
.param jc1end_r='jc1end*4'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='(max(1e-3,rendsh/multi/(wum-dwend))*tfacend)/2*(1+factmis)'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
rend1 n1 1  'rendo/2*(1+1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
r1 1 2  'ro/2*(3-1/(1+jc1_r1*v(1,2)*v(1,2)))'
r2 2 3  'ro*2/2*(3-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r3 3 4  'ro*2/2*(3-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r4 4 5  'ro*2/2*(3-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r5 5 6  'ro*2/2*(3-1/(1+jc1_r2*v(5,6)*v(5,6)))'
r6 6 7  'ro/2*(3-1/(1+jc1_r1*v(6,7)*v(6,7)))'
rend2 7 n2  'rendo/2*(1+1/(1+jc1end_r*v(7,n2)*v(7,n2)))'
d1 body 2 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
d2 body 3 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d3 body 4 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d4 body 5 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d5 body 6 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
.ends rnodwo_m
.subckt rpodwo_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00235891089108911*geo_fac*par_disres*mismatchflag'
.param rsh='r_rpodwo_m'     rendsh='2*rend_rpodwo_m*1e6'
.param dw_etch='0-0.0000000792*(pwr(0.545454545454545,x_dxw_rpodwo_m)-1)'
.param dw_emp='6.4000e-009'     dw_empend='2.2000e-008'
.param dl_etch='0+dxl_rpodwo_m'     dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'     dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=0.000045
.param jc1_w=0.000035     jc1_n=0.001
.param jc1end_0=0     jc1end_w=0
.param tc1_0=0.00105     tc1_w=9.088425e-07
.param tc2_0=1.0e-06     tc2_w=0
.param tc1end_0=0     tc1end_w=0
.param tc2end_0=0     tc2end_w=0
.param jct_0=0.00025     jct_w=0.0002
.param jct_n=0     jctend_0=0
.param jctend_w=0     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'     tc1='tc1_0 + tc1_w * min(wum, 5)'
.param tc2='tc2_0 + tc2_w * min(wum, 5)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 5)'
.param tc2end='tc2end_0 + tc2end_w * min(wum, 5)'
.param jct='jct_0 + jct_w * min(wum, 5) + jct_n * min(nsqr, 8)'
.param jctend='jctend_0 + jctend_w * min(wum, 5)'
.param jc1='(jc1_0 + jc1_w * min(wum, 5) + jc1_n * min(nsqr, 8) + jct * delta_t) / (lum-dl) / (lum-dl)'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param jc1end='max(0, (jc1end_0 + jc1end_w * min(wum, 5) + jctend * delta_t))'
.param jc1end_r='jc1end*4'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='(max(1e-3,rendsh/multi/(wum-dwend))*tfacend)/2*(1+factmis)'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
rend1 n1 1  'rendo/2*(3-1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
r1 1 2  'max(min(ro*(1+jc1_r1*v(1,2)*v(1,2)),ro*1.5),ro/2)'
r2 2 3  'max(min(ro*2*(1+jc1_r2*v(2,3)*v(2,3)),ro*3),ro)'
r3 3 4  'max(min(ro*2*(1+jc1_r2*v(3,4)*v(3,4)),ro*3),ro)'
r4 4 5  'max(min(ro*2*(1+jc1_r2*v(4,5)*v(4,5)),ro*3),ro)'
r5 5 6  'max(min(ro*2*(1+jc1_r2*v(5,6)*v(5,6)),ro*3),ro)'
r6 6 7  'max(min(ro*(1+jc1_r1*v(6,7)*v(6,7)),ro*1.5),ro/2)'
rend2 7 n2  'rendo/2*(3-1/(1+jc1end_r*v(7,n2)*v(7,n2)))'
d1 2 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
d2 3 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d3 4 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d4 5 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d5 6 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
.ends rpodwo_m
.subckt rnpolywo_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.025601414427157*geo_fac*par_disres*mismatchflag'
.param rsh='r_rnpolywo_m'     rendsh='2*rend_rnpolywo_m*1e6'
.param dw_etch='0-7.87500000000000e-008*(pwr(5.55555555555556e-001,x_dxw_rnpolywo_m)-1)'
.param dw_emp='1.8900e-008'     dw_empend='1.3800e-008'
.param dl_etch='0+dxl_rnpolywo_m'     dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'     dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=0.663686239758104
.param jc1_w=-0.0750065757208787     jc1_n=-0.000294462460888612
.param jc1end_0=13.3453193555066     jc1end_w=-0.175805407098847
.param tc1_0=0.000252907549762029     tc1_w=-1.09347086421216e-05
.param tc2_0=2.58388768423619e-07     tc2_w=-9.26075190896555e-10
.param tc1end_0=0.001764527883853     tc1end_w=-3.33638564578951e-06
.param tc2end_0=1.49538778703392e-07     tc2end_w=-3.81597136350383e-10
.param jct_0=0.000652309891571054     jct_w=-6.66283264583629e-05
.param jct_n=1.30784571473053e-07     jctend_0=-0.195545638318679
.param jctend_w=-0.122934918258964     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w / min(wum, 25)'
.param tc2='tc2_0 + tc2_w / min(wum, 25)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 25)'
.param tc2end='tc2end_0 + tc2end_w * min(wum, 25)'
.param jct='jct_0 + jct_w / min(wum, 25) + jct_n * min(nsqr, 150)'
.param jctend='jctend_0 + jctend_w * min(wum, 25)'
.param jc1='max(0, (jc1_0 + jc1_w / min(wum, 25) + jc1_n * min(nsqr, 150) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param jc1end='max(0, (jc1end_0 + jc1end_w / min(wum, 25) + jctend * delta_t))'
.param jc1end_r='jc1end*4'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='(max(1e-3,rendsh/multi/(wum-dwend))*tfacend)/2*(1+factmis)'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
.param ca=ca_pofox_r     cf=cf_polfox_r
.param af_rnpolywo_m=2
.param ef_rnpolywo_m=0.95
.param wf_rnpolywo_m=1
.param lf_rnpolywo_m=1
.param m_modfac='multi/(pwr(abs(multi),af_rnpolywo_m))'
.param a1_rnpolywo_m=4.25e-23
.param b1_rnpolywo_m=-1.7e-23
.param c1_rnpolywo_m=4.5e-23
.param kf_rnpolywo_m='(a1_rnpolywo_m*(abs(rnoiseflag_disres)+rnoiseflag_disres)+b1_rnpolywo_m*(abs(rnoiseflag_disres)-rnoiseflag_disres)+c1_rnpolywo_m)*m_modfac'
.model rnpoly1 r l='(lum-dl)*1e-6/10' w='(wum-dw)*1e-6' kf='kf_rnpolywo_m' af=af_rnpolywo_m ef=ef_rnpolywo_m wf=wf_rnpolywo_m lf=lf_rnpolywo_m
.model rnpoly2 r l='(lum-dl)*1e-6/5' w='(wum-dw)*1e-6' kf='kf_rnpolywo_m' af=af_rnpolywo_m ef=ef_rnpolywo_m wf=wf_rnpolywo_m lf=lf_rnpolywo_m
rend1 n1 1  'rendo/2*(3-1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
r1 1 2 rnpoly1 'ro/2*(3-1/(1+jc1_r1*v(1,2)*v(1,2)))'
r2 2 3 rnpoly2 'ro*2/2*(3-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r3 3 4 rnpoly2 'ro*2/2*(3-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r4 4 5 rnpoly2 'ro*2/2*(3-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r5 5 6 rnpoly2 'ro*2/2*(3-1/(1+jc1_r2*v(5,6)*v(5,6)))'
r6 6 7 rnpoly1 'ro/2*(3-1/(1+jc1_r1*v(6,7)*v(6,7)))'
rend2 7 n2  'rendo/2*(3-1/(1+jc1end_r*v(7,n2)*v(7,n2)))'
c1 body 2  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c2 body 3  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c3 body 4  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c4 body 5  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c5 body 6  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
.ends rnpolywo_m
.subckt rppolywo_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00545608203677511*geo_fac*par_disres*mismatchflag'
.param rsh='r_rppolywo_m'     rendsh='2*rend_rppolywo_m*1e6'
.param dw_etch='0-8.26333333333333e-008*(pwr(5.52238805970149e-001,x_dxw_rppolywo_m)-1)'
.param dw_emp='6.7280e-009'     dw_empend='-1.4670e-008'
.param dl_etch='0+dxl_rppolywo_m'     dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'     dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=0.0896111099341527
.param jc1_w=-0.00499080558384016     jc1_n=2.5374e-05
.param jc1end_0=6207.32004031375     jc1end_w=-1815.9
.param tc1_0=-0.000303589647270582     tc1_w=-1.12094842256059e-05
.param tc2_0=6.71216206685052e-07     tc2_w=2.2469040636621e-08
.param tc1end_0=-0.00113690867389968     tc1end_w=-0.000169845598239599
.param tc2end_0=1.3567176099377e-06     tc2end_w=-3.7427e-07
.param jct_0=-0.000412166544758672     jct_w=4.33890275487333e-05
.param jct_n=-1.9569e-09     jctend_0=-3.79298912034233
.param jctend_w=12.8609803922519     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w / min(wum, 25)'
.param tc2='tc2_0 + tc2_w / min(wum, 25)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 25)'
.param tc2end='tc2end_0 + tc2end_w * min(wum, 25)'
.param jct='jct_0 + jct_w / min(wum, 25) + jct_n * min(nsqr, 150)'
.param jctend='jctend_0 + jctend_w * min(wum, 25)'
.param jc1='max(0, (jc1_0 + jc1_w / min(wum, 25) + jc1_n * min(nsqr, 150) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param jc1end='max(0, (jc1end_0 + jc1end_w * min(wum, 25) + jctend * delta_t))'
.param jc1end_r='jc1end*4'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='(max(1e-3,rendsh/multi/(wum-dwend))*tfacend)/2*(1+factmis)'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
.param ca=ca_pofox_r     cf=cf_polfox_r
.param af_rppolywo_m=2
.param ef_rppolywo_m=0.95
.param wf_rppolywo_m=1
.param lf_rppolywo_m=1
.param m_modfac='multi/(pwr(abs(multi),af_rppolywo_m))'
.param a1_rppolywo_m=8.5e-23
.param b1_rppolywo_m=-3.1e-23
.param c1_rppolywo_m=1e-22
.param kf_rppolywo_m='(a1_rppolywo_m*(abs(rnoiseflag_disres)+rnoiseflag_disres)+b1_rppolywo_m*(abs(rnoiseflag_disres)-rnoiseflag_disres)+c1_rppolywo_m)*m_modfac'
.model rppoly1 r l='(lum-dl)*1e-6/10' w='(wum-dw)*1e-6' kf='kf_rppolywo_m' af=af_rppolywo_m ef=ef_rppolywo_m wf=wf_rppolywo_m lf=lf_rppolywo_m
.model rppoly2 r l='(lum-dl)*1e-6/5' w='(wum-dw)*1e-6' kf='kf_rppolywo_m' af=af_rppolywo_m ef=ef_rppolywo_m wf=wf_rppolywo_m lf=lf_rppolywo_m
rend1 n1 1  'rendo/2*(3-1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
r1 1 2 rppoly1 'ro/2*(1+1/(1+jc1_r1*v(1,2)*v(1,2)))'
r2 2 3 rppoly2 'ro*2/2*(1+1/(1+jc1_r2*v(2,3)*v(2,3)))'
r3 3 4 rppoly2 'ro*2/2*(1+1/(1+jc1_r2*v(3,4)*v(3,4)))'
r4 4 5 rppoly2 'ro*2/2*(1+1/(1+jc1_r2*v(4,5)*v(4,5)))'
r5 5 6 rppoly2 'ro*2/2*(1+1/(1+jc1_r2*v(5,6)*v(5,6)))'
r6 6 7 rppoly1 'ro/2*(1+1/(1+jc1_r1*v(6,7)*v(6,7)))'
rend2 7 n2  'rendo/2*(3-1/(1+jc1end_r*v(7,n2)*v(7,n2)))'
c1 body 2  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c2 body 3  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c3 body 4  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c4 body 5  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c5 body 6  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
.ends rppolywo_m
.subckt rnodl_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00388246110325318*geo_fac*par_disres*mismatchflag'
.param rsh='r_rnodl_m'
.param dw_etch='0-1.51144067796610e-008*(pwr(abs(+4.24390243902439e-001),x_dxw_rnodl_m)-1)'
.param dw_emp='-1.7500e-008'     dl_etch='0+dxl_rnodl_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=2.29716374936608
.param jc1_w=0.966849672886205     jc1_n=-0.00186855903400384
.param tc1_0=0.00163137853390732     tc1_w=-2.06701587598843e-06
.param tc2_0=4.59142442126849e-10     tc2_w=-2.20926894845178e-09
.param jct_0=-0.00367376044027522     jct_w=0.000927708589609838
.param jct_n=6.00355804266836e-07     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
r1 n1 1  'ro/2*(3-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2/2*(3-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2/2*(3-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2/2*(3-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2/2*(3-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro/2*(3-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
d1 body 1 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
d2 body 2 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d3 body 3 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d4 body 4 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d5 body 5 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
.ends rnodl_m
.subckt rnods_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00388246110325318*geo_fac*par_disres*mismatchflag'
.param rsh='r_rnods_m'
.param dw_etch='0-1.51144067796610e-008*(pwr(abs(+4.24390243902439e-001),x_dxw_rnods_m)-1)'
.param dw_emp='-1.7500e-008'     dl_etch='0+dxl_rnods_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=2.29716374936608
.param jc1_w=0.966849672886205     jc1_n=-0.00186855903400384
.param tc1_0=0.00163137853390732     tc1_w=-2.06701587598843e-06
.param tc2_0=4.59142442126849e-10     tc2_w=-2.20926894845178e-09
.param jct_0=-0.00367376044027522     jct_w=0.000927708589609838
.param jct_n=6.00355804266836e-07     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
r1 n1 1  'ro/2*(3-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2/2*(3-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2/2*(3-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2/2*(3-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2/2*(3-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro/2*(3-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
d1 body 1 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
d2 body 2 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d3 body 3 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d4 body 4 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d5 body 5 ndio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
.ends rnods_m
.subckt rpodl_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00646096181046676*geo_fac*par_disres*mismatchflag'
.param rsh='r_rpodl_m'
.param dw_etch='0-7.64533333333333e-009*(pwr(abs(+3.85245901639344e-001),x_dxw_rpodl_m)-1)'
.param dw_emp='-1.8000e-008'     dl_etch='0+dxl_rpodl_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=2.43769875284375
.param jc1_w=0.958671839463289     jc1_n=-0.000527375464451339
.param tc1_0=0.00205     tc1_w=-7e-04
.param tc2_0=-7.71968996056192e-08     tc2_w=-5.17108135853353e-09
.param jct_0=-0.00402689298858613     jct_w=0.000741523846651567
.param jct_n=-3.97127786494667e-06     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 0.5)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param drsh=0     rshh=0.21
.param rshn=1     ww=0
.param wwn=1     deltar='drsh+rshh/pwr(wum,rshn)'
.param deltaw='dw+ww/pwr(wum,wwn)'     reff='(rsh-deltar)'
.param ro='(reff/multi*(lum-dl)/(wum-deltaw)*tfac)/10*(1+factmis)'
r1 n1 1  'ro/2*(3-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2/2*(3-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2/2*(3-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2/2*(3-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2/2*(3-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro/2*(3-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
d1 1 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
d2 2 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d3 3 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d4 4 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d5 5 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
.ends rpodl_m
.subckt rpods_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00646096181046676*geo_fac*par_disres*mismatchflag'
.param rsh='r_rpods_m'
.param dw_etch='0-7.64533333333333e-009*(pwr(abs(+3.85245901639344e-001),x_dxw_rpods_m)-1)'
.param dw_emp='-1.8000e-008'     dl_etch='0+dxl_rpods_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=2.43769875284375
.param jc1_w=0.958671839463289     jc1_n=-0.000527375464451339
.param tc1_0=0.00205     tc1_w=-7e-04
.param tc2_0=-7.71968996056192e-08     tc2_w=-5.17108135853353e-09
.param jct_0=-0.00402689298858613     jct_w=0.000741523846651567
.param jct_n=-3.97127786494667e-06     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 0.5)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param drsh=0     rshh=0.21
.param rshn=1     ww=0
.param wwn=1     deltar='drsh+rshh/pwr(wum,rshn)'
.param deltaw='dw+ww/pwr(wum,wwn)'     reff='(rsh-deltar)'
.param ro='(reff/multi*(lum-dl)/(wum-deltaw)*tfac)/10*(1+factmis)'
r1 n1 1  'ro/2*(3-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2/2*(3-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2/2*(3-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2/2*(3-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2/2*(3-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro/2*(3-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
d1 1 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
d2 2 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d3 3 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d4 4 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*(2.0*(lr-dl/scale*1e-6)/5.0)'
d5 5 body pdio  area='multi*((wr-dw/scale*1e-6)*(lr-dl/scale*1e-6)/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*(lr-dl/scale*1e-6)/5.0)'
.ends rpods_m
.subckt rnpolyl_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00617892503536068*geo_fac*par_disres*mismatchflag'
.param rsh='r_rnpolyl_m'
.param dw_etch='0-6.52202838557067e-009*(pwr(abs(+4.25025501530092e-001),x_dxw_rnpolyl_m)-1)'
.param dw_emp='2.6400e-009'     dl_etch='0+dxl_rnpolyl_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=6.5
.param jc1_w=5.9     jc1_n=-7e-3
.param tc1_0=0.00160199933242697     tc1_w=-1.2104e-05
.param tc2_0=1.1174e-07     tc2_w=2.5013e-08
.param jct_0=-0.0185506445636512     jct_w=-0.0334478918733522
.param jct_n=3.1771e-05     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 1) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 3) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
.param ca=ca_pofox     cf=cf_polfox
r1 n1 1  'ro*(2-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2*(2-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2*(2-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2*(2-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2*(2-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro*(2-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
c1 body 1  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c2 body 2  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c3 body 3  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c4 body 4  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c5 body 5  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
.ends rnpolyl_m
.subckt rnpolys_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00617892503536068*geo_fac*par_disres*mismatchflag'
.param rsh='r_rnpolys_m'
.param dw_etch='0-6.52202838557067e-009*(pwr(abs(+4.25025501530092e-001),x_dxw_rnpolys_m)-1)'
.param dw_emp='2.6400e-009'     dl_etch='0+dxl_rnpolys_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=6.5
.param jc1_w=5.9     jc1_n=-7e-3
.param tc1_0=0.00160199933242697     tc1_w=-1.2104e-05
.param tc2_0=1.1174e-07     tc2_w=2.5013e-08
.param jct_0=-0.0185506445636512     jct_w=-0.0334478918733522
.param jct_n=3.1771e-05     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 1) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 3) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
.param ca=ca_pofox     cf=cf_posfox
r1 n1 1  'ro*(2-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2*(2-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2*(2-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2*(2-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2*(2-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro*(2-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
c1 body 1  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c2 body 2  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c3 body 3  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c4 body 4  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c5 body 5  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
.ends rnpolys_m
.subckt rppolyl_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00706718528995757*geo_fac*par_disres*mismatchflag'
.param rsh='r_rppolyl_m'
.param dw_etch='0-7.92704402515723e-009*(pwr(abs(+4.19708029197080e-001),x_dxw_rppolyl_m)-1)'
.param dw_emp='-5.1000e-009'     dl_etch='0+dxl_rppolyl_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=9.5
.param jc1_w=5.81508402119467     jc1_n=-0.00923267200801938
.param tc1_0=0.00194430976641791     tc1_w=-5.15825498692349e-05
.param tc2_0=1.6539e-07     tc2_w=1.2637e-08
.param jct_0=-0.0460444710839901     jct_w=-1.8e-2
.param jct_n=4.3569e-05     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'     tc1='tc1_0 + tc1_w * min(wum, 5)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 2) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 4) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
.param ca=ca_pofox     cf=cf_polfox
r1 n1 1  'ro*(2-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2*(2-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2*(2-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2*(2-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2*(2-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro*(2-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
c1 body 1  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c2 body 2  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c3 body 3  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c4 body 4  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c5 body 5  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
.ends rppolyl_m
.subckt rppolys_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres' mismatchflag='mismatchflag_disres'
.param geo_fac='1/sqrt(multi*lr*scale*wr*scale*1e12)'
.param factmis='0.00706718528995757*geo_fac*par_disres*mismatchflag'
.param rsh='r_rppolys_m'
.param dw_etch='0-7.92704402515723e-009*(pwr(abs(+4.19708029197080e-001),x_dxw_rppolys_m)-1)'
.param dw_emp='-5.1000e-009'     dl_etch='0+dxl_rppolys_m'
.param dxl_r='0.0000e+000'     dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'     jc1_0=9.5
.param jc1_w=5.81508402119467     jc1_n=-0.00923267200801938
.param tc1_0=0.00194430976641791     tc1_w=-5.15825498692349e-05
.param tc2_0=1.6539e-07     tc2_w=1.2637e-08
.param jct_0=-0.0460444710839901     jct_w=-1.8e-2
.param jct_n=4.3569e-05     delta_t='temper - 25'
.param lum='lr*scale*1e6'     wum='wr*scale*1e6'
.param nsqr='lr/wr'     tc1='tc1_0 + tc1_w * min(wum, 5)'
.param tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 2) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 4) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r1='jc1*100'     jc1_r2='jc1*25'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='(max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac)/10*(1+factmis)'
.param ca=ca_pofox     cf=cf_posfox
r1 n1 1  'ro*(2-1/(1+jc1_r1*v(n1,1)*v(n1,1)))'
r2 1 2  'ro*2*(2-1/(1+jc1_r2*v(1,2)*v(1,2)))'
r3 2 3  'ro*2*(2-1/(1+jc1_r2*v(2,3)*v(2,3)))'
r4 3 4  'ro*2*(2-1/(1+jc1_r2*v(3,4)*v(3,4)))'
r5 4 5  'ro*2*(2-1/(1+jc1_r2*v(4,5)*v(4,5)))'
r6 5 n2  'ro*(2-1/(1+jc1_r1*v(5,n2)*v(5,n2)))'
c1 body 1  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c2 body 2  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c3 body 3  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c4 body 4  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
c5 body 5  'multi*(ca*((wr*scale)*lr*scale/5.0)*1e12+2*cf*lr*scale/5.0*1e6)'
.ends rppolys_m
.subckt rnwod_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres'
.param rsh=r_rnwod_m     dw=0.135u
.param pt='temper'
.param pvc1='(1.993e-08/(max(wr*scale*1e6,1.8))+1.259e-09)*(min(lr*scale*1e6,50))+(-5.381e-08/(max(wr*scale*1e6,1.8))+6.448e-08)'
.param pvc1_r1='pvc1*10'     pvc1_r2='pvc1*5'
.param pvc2=0     pvc2_r1='pvc2*100'
.param pvc2_r2='pvc2*25'     ptc1=1.951e-03
.param ptc2=8.526e-06
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
.param rmain='(rsh/multi*lr*scale/(wr*scale-dw)*tfac)/10'
.param rend='rend_rnwod_m'
rend1 n1 1  'rend/multi/(wr*scale+0.5u)'
r1 1 2  'max(min(rmain*(1+pvc1_r1*(abs(v(1,2))/lr/scale)+pvc2_r1*(v(1,2)/lr/scale)*(v(1,2)/lr/scale)),rmain*1.5),rmain/2)'
r2 2 3  'max(min(rmain*2*(1+pvc1_r2*(abs(v(2,3))/lr/scale)+pvc2_r2*(v(2,3)/lr/scale)*(v(2,3)/lr/scale)),rmain*3),rmain)'
r3 3 4  'max(min(rmain*2*(1+pvc1_r2*(abs(v(3,4))/lr/scale)+pvc2_r2*(v(3,4)/lr/scale)*(v(3,4)/lr/scale)),rmain*3),rmain)'
r4 4 5  'max(min(rmain*2*(1+pvc1_r2*(abs(v(4,5))/lr/scale)+pvc2_r2*(v(4,5)/lr/scale)*(v(4,5)/lr/scale)),rmain*3),rmain)'
r5 5 6  'max(min(rmain*2*(1+pvc1_r2*(abs(v(5,6))/lr/scale)+pvc2_r2*(v(5,6)/lr/scale)*(v(5,6)/lr/scale)),rmain*3),rmain)'
r6 6 7  'max(min(rmain*(1+pvc1_r1*(abs(v(6,7))/lr/scale)+pvc2_r1*(v(6,7)/lr/scale)*(v(6,7)/lr/scale)),rmain*1.5),rmain/2)'
rend2 7 n2  'rend/multi/(wr*scale+0.5u)'
d1 body 2 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*lr/5.0)'
d2 body 3 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*2.0*lr/5.0'
d3 body 4 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*2.0*lr/5.0'
d4 body 5 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*2.0*lr/5.0'
d5 body 6 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*lr/5.0)'
.ends rnwod_m
.subckt rnwsti_m n1 n2 body lr=length wr=width multi=1 scale='scale_disres'
.param rsh=r_rnwsti_m     dw=3.68e-7
.param pt='temper'
.param pvc1='(3.369e-08/(max(wr*scale*1e6,1.8))+8.881e-10)*(min(lr*scale*1e6,50))+(-1.492e-07/(max(wr*scale*1e6,1.8))+1.8e-07)'
.param pvc1_r1='pvc1*10'     pvc1_r2='pvc1*5'
.param pvc2=0     pvc2_r1='pvc2*100'
.param pvc2_r2='pvc2*25'     ptc1=2.806e-03
.param ptc2=8.932e-06
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
.param rmain='(rsh/multi*lr*scale/(wr*scale-dw)*tfac)/10'
.param rend='rend_rnwsti_m'
rend1 n1 1  'rend/multi/(wr*scale)'
r1 1 2  'max(min(rmain*(1+pvc1_r1*(abs(v(1,2))/lr/scale)+pvc2_r1*(v(1,2)/lr/scale)*(v(1,2)/lr/scale)),rmain*1.5),rmain/2)'
r2 2 3  'max(min(rmain*2*(1+pvc1_r2*(abs(v(2,3))/lr/scale)+pvc2_r2*(v(2,3)/lr/scale)*(v(2,3)/lr/scale)),rmain*3),rmain)'
r3 3 4  'max(min(rmain*2*(1+pvc1_r2*(abs(v(3,4))/lr/scale)+pvc2_r2*(v(3,4)/lr/scale)*(v(3,4)/lr/scale)),rmain*3),rmain)'
r4 4 5  'max(min(rmain*2*(1+pvc1_r2*(abs(v(4,5))/lr/scale)+pvc2_r2*(v(4,5)/lr/scale)*(v(4,5)/lr/scale)),rmain*3),rmain)'
r5 5 6  'max(min(rmain*2*(1+pvc1_r2*(abs(v(5,6))/lr/scale)+pvc2_r2*(v(5,6)/lr/scale)*(v(5,6)/lr/scale)),rmain*3),rmain)'
r6 6 7  'max(min(rmain*(1+pvc1_r1*(abs(v(6,7))/lr/scale)+pvc2_r1*(v(6,7)/lr/scale)*(v(6,7)/lr/scale)),rmain*1.5),rmain/2)'
rend2 7 n2  'rend/multi/(wr*scale)'
d1 body 2 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*lr/5.0)'
d2 body 3 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*2.0*lr/5.0'
d3 body 4 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*2.0*lr/5.0'
d4 body 5 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*2.0*lr/5.0'
d5 body 6 nwdio  area='multi*((wr-dw/scale*1e-6)*lr/5.0)' pj='multi*((wr-dw/scale*1e-6)+2.0*lr/5.0)'
.ends rnwsti_m
.param mismatchflag_res=1
.param scale_res=0.9
.param rnoiseflag_res=0
.param par_res=agauss(0,1,1) r_rnodwo=1.0930e+002       rend_rnodwo=9.5824e-006        x_dxw_rnodwo=0         dxl_rnodwo=0 r_rpodwo=3.1373e+002       rend_rpodwo=6.0000e-006        x_dxw_rpodwo=0         dxl_rpodwo=0 r_rnpolywo=1.4970e+002     rend_rnpolywo=7.5700e-006      x_dxw_rnpolywo=0     dxl_rnpolywo=0 r_rppolywo=8.7600e+002     rend_rppolywo=6.2372e-006      x_dxw_rppolywo=0     dxl_rppolywo=0 r_rnodl=1.8000e+001            dxl_rnodl=0       x_dxw_rnodl=0 r_rnods=1.8000e+001            dxl_rnods=0       x_dxw_rnods=0 r_rpodl=1.6700e+001            dxl_rpodl=0       x_dxw_rpodl=0 r_rpods=1.6700e+001            dxl_rpods=0       x_dxw_rpods=0 r_rnpolyl=1.6420e+001          dxl_rnpolyl=0     x_dxw_rnpolyl=0 r_rnpolys=1.6420e+001          dxl_rnpolys=0     x_dxw_rnpolys=0 r_rppolyl=1.4400e+001          dxl_rppolyl=0     x_dxw_rppolyl=0 r_rppolys=1.4400e+001          dxl_rppolys=0     x_dxw_rppolys=0 r_rnwod=385            rend_rnwod='170e-6' r_rnwsti=1169           rend_rnwsti='2.7e-4' r_rm1l=0.136             r_rm1s=0.308             r_rm1w=0.225 r_rm2l=0.13              r_rm2s=0.292             r_rm2w=0.21 r_rm3l=0.13              r_rm3s=0.292             r_rm3w=0.21 r_rm4l=0.13              r_rm4s=0.292             r_rm4w=0.21 r_rm5l=0.13              r_rm5s=0.292             r_rm5w=0.21 r_rm6l=0.13              r_rm6s=0.292             r_rm6w=0.21 r_rm7l=0.13              r_rm7s=0.292             r_rm7w=0.21 r_rm8l=0.13              r_rm8s=0.292             r_rm8w=0.21 r_rm9l=0.0221            r_rm9s=0.0218            r_rm9w=0.0229 r_rm10l=0.0221            r_rm10s=0.0218            r_rm10w=0.0229 r_rm11=0.0183            r_rmxl=0.13              r_rmxs=0.292 r_rmxw=0.21              r_rmyl=0.0683            r_rmys=0.1002 r_rmyw=0.0827            r_rmytl=0.0599            r_rmyts=0.095 r_rmytw=0.0772            r_rmzl=0.0221            r_rmzs=0.0218 r_rmzw=0.0229            r_rmrl=0.0167            r_rmrs=0.0165 r_rmrw=0.0175
.subckt rnodwo n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00198323903818953*geo_fac*par_res*mismatchflag'
.param rsh='r_rnodwo'  rendsh='2*rend_rnodwo*1e6'
.param dw_etch='0-9.25714285714286e-08*(pwr(0.5625,x_dxw_rnodwo)-1)'   dw_emp='1.5370e-009'    dw_empend='-5.2360e-008'
.param dl_etch='0+dxl_rnodwo'      dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'  dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=0.411133860400214  jc1_w=0.0577271204979308  jc1_n=-0.00313
.param jc1end_0=-1.13929  jc1end_w=40.82881
.param tc1_0=0.0014342814911298  tc1_w=-2.24331695355166e-07
.param tc2_0=7.54746914856436e-07  tc2_w=-2.0217e-09
.param tc1end_0=0.00135719397917256  tc1end_w=2.1275e-05
.param tc2end_0=3.37552662511097e-07  tc2end_w=-1.481e-08
.param jct_0=-0.00027337  jct_w=0.00019370448410292  jct_n=-3.8271e-06
.param jctend_0=-0.0487  jctend_w=0.0962829566646918
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 25)'   tc2='tc2_0 + tc2_w * min(wum, 25)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 25)'   tc2end='tc2end_0 + tc2end_w * min(wum, 25)'
.param jct='jct_0 + jct_w * min(wum, 25) + jct_n * min(nsqr, 150)'
.param jctend='jctend_0 + jctend_w * min(wum, 25)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 25) + jc1_n * min(nsqr, 150) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param jc1end='max(0, (jc1end_0 + jc1end_w * min(wum, 25) + jctend * delta_t))'
.param jc1end_r='jc1end'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='max(1e-3,rendsh/multi/(wum-dwend))*tfacend*(1+factmis)'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rend n1 1 'rendo/2*(1+1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
rmain 1 n2 'ro/2*(3-1/(1+jc1_r*v(1,n2)*v(1,n2)))'
.ends rnodwo
.subckt rpodwo n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00235891089108911*geo_fac*par_res*mismatchflag'
.param rsh='r_rpodwo'  rendsh='2*rend_rpodwo*1e6'
.param dw_etch='0-0.0000000792*(pwr(0.545454545454545,x_dxw_rpodwo)-1)'   dw_emp='6.4000e-009'     dw_empend='2.2000e-008'
.param dl_etch='0+dxl_rpodwo'      dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'  dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=0.000045  jc1_w=0.000035   jc1_n=0.001
.param jc1end_0=0 jc1end_w=0
.param tc1_0=0.00105  tc1_w=9.088425e-07
.param tc2_0=1.0e-06  tc2_w=0
.param tc1end_0=0  tc1end_w=0
.param tc2end_0=0  tc2end_w=0
.param jct_0=0.00025  jct_w=0.0002 jct_n=0
.param jctend_0=0  jctend_w=0
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 5)'   tc2='tc2_0 + tc2_w * min(wum, 5)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 5)'   tc2end='tc2end_0 + tc2end_w * min(wum, 5)'
.param jct='jct_0 + jct_w * min(wum, 5) + jct_n * min(nsqr, 8)'
.param jctend='jctend_0 + jctend_w * min(wum, 5)'
.param jc1='(jc1_0 + jc1_w * min(wum, 5) + jc1_n * min(nsqr, 8) + jct * delta_t) / (lum-dl) / (lum-dl)'
.param jc1_r='jc1'
.param jc1end='max(0, (jc1end_0 + jc1end_w * min(wum, 5) + jctend * delta_t))'
.param jc1end_r='jc1end'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='max(1e-3,rendsh/multi/(wum-dwend))*tfacend*(1+factmis)'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rend n1 1 'rendo/2*(3-1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
rmain 1 n2 'max(min(ro*(1+jc1_r*v(1,n2)*v(1,n2)), ro*1.5), ro/2)'
.ends rpodwo
.subckt rnpolywo n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.025601414427157*geo_fac*par_res*mismatchflag'
.param rsh='r_rnpolywo'  rendsh='2*rend_rnpolywo*1e6'
.param dw_etch='0-7.87500000000000e-008*(pwr(5.55555555555556e-001,x_dxw_rnpolywo)-1)'   dw_emp='1.8900e-008'    dw_empend='1.3800e-008'
.param dl_etch='0+dxl_rnpolywo'     dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'  dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=0.663686239758104  jc1_w=-0.0750065757208787  jc1_n=-0.000294462460888612
.param jc1end_0=13.3453193555066  jc1end_w=-0.175805407098847
.param tc1_0=0.000252907549762029  tc1_w=-1.09347086421216e-05
.param tc2_0=2.58388768423619e-07  tc2_w=-9.26075190896555e-10
.param tc1end_0=0.001764527883853  tc1end_w=-3.33638564578951e-06
.param tc2end_0=1.49538778703392e-07  tc2end_w=-3.81597136350383e-10
.param jct_0=0.000652309891571054  jct_w=-6.66283264583629e-05  jct_n=1.30784571473053e-07
.param jctend_0=-0.195545638318679  jctend_w=-0.122934918258964
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w / min(wum, 25)'   tc2='tc2_0 + tc2_w / min(wum, 25)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 25)'   tc2end='tc2end_0 + tc2end_w * min(wum, 25)'
.param jct='jct_0 + jct_w / min(wum, 25) + jct_n * min(nsqr, 150)'
.param jctend='jctend_0 + jctend_w * min(wum, 25)'
.param jc1='max(0, (jc1_0 + jc1_w / min(wum, 25) + jc1_n * min(nsqr, 150) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param jc1end='max(0, (jc1end_0 + jc1end_w / min(wum, 25) + jctend * delta_t))'
.param jc1end_r='jc1end'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='max(1e-3,rendsh/multi/(wum-dwend))*tfacend*(1+factmis)'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
.param af_rnpolywo=2
.param ef_rnpolywo=0.95
.param wf_rnpolywo=1
.param lf_rnpolywo=1
.param m_modfac='multi/(pwr(abs(multi),af_rnpolywo))'
.param a1_rnpolywo=4.25e-23
.param b1_rnpolywo=-1.7e-23
.param c1_rnpolywo=4.5e-23
.param kf_rnpolywo='(a1_rnpolywo*(abs(rnoiseflag_res)+rnoiseflag_res)+b1_rnpolywo*(abs(rnoiseflag_res)-rnoiseflag_res)+c1_rnpolywo)*m_modfac'
rend n1 1 'rendo/2*(3-1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
rmain 1 n2 rnpoly 'ro/2*(3-1/(1+jc1_r*v(1,n2)*v(1,n2)))'
.model rnpoly r l='(lum-dl)*1e-6/1' w='(wum-dw)*1e-6' kf='kf_rnpolywo' af=af_rnpolywo ef=ef_rnpolywo wf=wf_rnpolywo lf=lf_rnpolywo
.ends rnpolywo
.subckt rppolywo n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00545608203677511*geo_fac*par_res*mismatchflag'
.param rsh='r_rppolywo'  rendsh='2*rend_rppolywo*1e6'
.param dw_etch='0-8.26333333333333e-008*(pwr(5.52238805970149e-001,x_dxw_rppolywo)-1)'    dw_emp='6.7280e-009'    dw_empend='-1.4670e-008'
.param dl_etch='0+dxl_rppolywo'       dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'  dwend='(dw_etch+dw_empend)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=0.0896111099341527  jc1_w=-0.00499080558384016  jc1_n=2.5374e-05
.param jc1end_0=6207.32004031375  jc1end_w=-1815.9
.param tc1_0=-0.000303589647270582  tc1_w=-1.12094842256059e-05
.param tc2_0=6.71216206685052e-07  tc2_w=2.2469040636621e-08
.param tc1end_0=-0.00113690867389968  tc1end_w=-0.000169845598239599
.param tc2end_0=1.3567176099377e-06  tc2end_w=-3.7427e-07
.param jct_0=-0.000412166544758672  jct_w=4.33890275487333e-05  jct_n=-1.9569e-09
.param jctend_0=-3.79298912034233  jctend_w=12.8609803922519
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w / min(wum, 25)'   tc2='tc2_0 + tc2_w / min(wum, 25)'
.param tc1end='tc1end_0 + tc1end_w * min(wum, 25)'   tc2end='tc2end_0 + tc2end_w * min(wum, 25)'
.param jct='jct_0 + jct_w / min(wum, 25) + jct_n * min(nsqr, 150)'
.param jctend='jctend_0 + jctend_w * min(wum, 25)'
.param jc1='max(0, (jc1_0 + jc1_w / min(wum, 25) + jc1_n * min(nsqr, 150) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param jc1end='max(0, (jc1end_0 + jc1end_w * min(wum, 25) + jctend * delta_t))'
.param jc1end_r='jc1end'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param tfacend='1 + tc1end * delta_t + tc2end * delta_t * delta_t'
.param rendo='max(1e-3,rendsh/multi/(wum-dwend))*tfacend*(1+factmis)'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
.param af_rppolywo=2
.param ef_rppolywo=0.95
.param wf_rppolywo=1
.param lf_rppolywo=1
.param m_modfac='multi/(pwr(abs(multi),af_rppolywo))'
.param a1_rppolywo=8.5e-23
.param b1_rppolywo=-3.1e-23
.param c1_rppolywo=1e-22
.param kf_rppolywo='(a1_rppolywo*(abs(rnoiseflag_res)+rnoiseflag_res)+b1_rppolywo*(abs(rnoiseflag_res)-rnoiseflag_res)+c1_rppolywo)*m_modfac'
rend n1 1 'rendo/2*(3-1/(1+jc1end_r*v(n1,1)*v(n1,1)))'
rmain 1 n2 rppoly 'ro/2*(1+1/(1+jc1_r*v(1,n2)*v(1,n2)))'
.model rppoly r l='(lum-dl)*1e-6/1' w='(wum-dw)*1e-6' kf='kf_rppolywo' af=af_rppolywo ef=ef_rppolywo wf=wf_rppolywo lf=lf_rppolywo
.ends rppolywo
.subckt rnodl n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00388246110325318*geo_fac*par_res*mismatchflag'
.param rsh='r_rnodl'
.param dw_etch='0-1.51144067796610e-008*(pwr(abs(+4.24390243902439e-001),x_dxw_rnodl)-1)'     dw_emp='-1.7500e-008'
.param dl_etch='0+dxl_rnodl'      dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=2.29716374936608  jc1_w=0.966849672886205  jc1_n=-0.00186855903400384
.param tc1_0=0.00163137853390732  tc1_w=-2.06701587598843e-06
.param tc2_0=4.59142442126849e-10  tc2_w=-2.20926894845178e-09
.param jct_0=-0.00367376044027522  jct_w=0.000927708589609838  jct_n=6.00355804266836e-07
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rmain n1 n2 'ro/2*(3-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rnodl
.subckt rnods n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00388246110325318*geo_fac*par_res*mismatchflag'
.param rsh='r_rnods'
.param dw_etch='0-1.51144067796610e-008*(pwr(abs(+4.24390243902439e-001),x_dxw_rnods)-1)'     dw_emp='-1.7500e-008'
.param dl_etch='0+dxl_rnods'      dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=2.29716374936608  jc1_w=0.966849672886205  jc1_n=-0.00186855903400384
.param tc1_0=0.00163137853390732  tc1_w=-2.06701587598843e-06
.param tc2_0=4.59142442126849e-10  tc2_w=-2.20926894845178e-09
.param jct_0=-0.00367376044027522  jct_w=0.000927708589609838  jct_n=6.00355804266836e-07
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rmain n1 n2 'ro/2*(3-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rnods
.subckt rpodl n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00646096181046676*geo_fac*par_res*mismatchflag'
.param rsh='r_rpodl'
.param dw_etch='0-7.64533333333333e-009*(pwr(abs(+3.85245901639344e-001),x_dxw_rpodl)-1)'          dw_emp='-1.8000e-008'
.param dl_etch='0+dxl_rpodl'            dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=2.43769875284375  jc1_w=0.958671839463289  jc1_n=-0.000527375464451339
.param tc1_0=0.00205  tc1_w=-7e-04
.param tc2_0=-7.71968996056192e-08  tc2_w=-5.17108135853353e-09
.param jct_0=-0.00402689298858613  jct_w=0.000741523846651567  jct_n=-3.97127786494667e-06
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 0.5)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param drsh=0    rshh=0.21    rshn=1
.param ww=0    wwn=1
.param deltar='drsh+rshh/pwr(wum,rshn)'
.param deltaw='dw+ww/pwr(wum,wwn)'
.param reff='(rsh-deltar)'
.param ro='reff/multi*(lum-dl)/(wum-deltaw)*tfac*(1+factmis)'
rmain n1 n2 'ro/2*(3-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rpodl
.subckt rpods n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00646096181046676*geo_fac*par_res*mismatchflag'
.param rsh='r_rpods'
.param dw_etch='0-7.64533333333333e-009*(pwr(abs(+3.85245901639344e-001),x_dxw_rpods)-1)'          dw_emp='-1.8000e-008'
.param dl_etch='0+dxl_rpods'            dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=2.43769875284375  jc1_w=0.958671839463289  jc1_n=-0.000527375464451339
.param tc1_0=0.00205  tc1_w=-7e-04
.param tc2_0=-7.71968996056192e-08  tc2_w=-5.17108135853353e-09
.param jct_0=-0.00402689298858613  jct_w=0.000741523846651567  jct_n=-3.97127786494667e-06
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 0.5)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 10) + jct_n * min(nsqr, 727.272727272727)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 10) + jc1_n * min(nsqr, 727.272727272727) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param drsh=0    rshh=0.21    rshn=1
.param ww=0    wwn=1
.param deltar='drsh+rshh/pwr(wum,rshn)'
.param deltaw='dw+ww/pwr(wum,wwn)'
.param reff='(rsh-deltar)'
.param ro='reff/multi*(lum-dl)/(wum-deltaw)*tfac*(1+factmis)'
rmain n1 n2 'ro/2*(3-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rpods
.subckt rnpolyl n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00617892503536068*geo_fac*par_res*mismatchflag'
.param rsh='r_rnpolyl'
.param dw_etch='0-6.52202838557067e-009*(pwr(abs(+4.25025501530092e-001),x_dxw_rnpolyl)-1)'       dw_emp='2.6400e-009'
.param dl_etch='0+dxl_rnpolyl'           dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=6.5  jc1_w=5.9  jc1_n=-7e-3
.param tc1_0=0.00160199933242697  tc1_w=-1.2104e-05
.param tc2_0=1.1174e-07  tc2_w=2.5013e-08
.param jct_0=-0.0185506445636512  jct_w=-0.0334478918733522  jct_n=3.1771e-05
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 1) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 3) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rmain n1 n2 'ro*(2-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rnpolyl
.subckt rnpolys n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00617892503536068*geo_fac*par_res*mismatchflag'
.param rsh='r_rnpolys'
.param dw_etch='0-6.52202838557067e-009*(pwr(abs(+4.25025501530092e-001),x_dxw_rnpolys)-1)'       dw_emp='2.6400e-009'
.param dl_etch='0+dxl_rnpolys'           dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=6.5  jc1_w=5.9  jc1_n=-7e-3
.param tc1_0=0.00160199933242697  tc1_w=-1.2104e-05
.param tc2_0=1.1174e-07  tc2_w=2.5013e-08
.param jct_0=-0.0185506445636512  jct_w=-0.0334478918733522  jct_n=3.1771e-05
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 10)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 1) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 3) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rmain n1 n2 'ro*(2-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rnpolys
.subckt rppolyl n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00706718528995757*geo_fac*par_res*mismatchflag'
.param rsh='r_rppolyl'
.param dw_etch='0-7.92704402515723e-009*(pwr(abs(+4.19708029197080e-001),x_dxw_rppolyl)-1)'   dw_emp='-5.1000e-009'
.param dl_etch='0+dxl_rppolyl'        dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=9.5  jc1_w=5.81508402119467  jc1_n=-0.00923267200801938
.param tc1_0=0.00194430976641791  tc1_w=-5.15825498692349e-05
.param tc2_0=1.6539e-07  tc2_w=1.2637e-08
.param jct_0=-0.0460444710839901  jct_w=-1.8e-2 jct_n=4.3569e-05
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 5)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 2) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 4) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rmain n1 n2 'ro*(2-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rppolyl
.subckt rppolys n1 n2 l=length w=width scale='scale_res' multi=1 mismatchflag='mismatchflag_res'
.param geo_fac='1/sqrt(multi*l*scale*w*scale*1e12)'
.param factmis='0.00706718528995757*geo_fac*par_res*mismatchflag'
.param rsh='r_rppolys'
.param dw_etch='0-7.92704402515723e-009*(pwr(abs(+4.19708029197080e-001),x_dxw_rppolys)-1)'   dw_emp='-5.1000e-009'
.param dl_etch='0+dxl_rppolys'        dxl_r='0.0000e+000'
.param dw='(dw_etch+dw_emp)*1e6'
.param dl='(dl_etch+dxl_r)*1e6'
.param jc1_0=9.5  jc1_w=5.81508402119467  jc1_n=-0.00923267200801938
.param tc1_0=0.00194430976641791  tc1_w=-5.15825498692349e-05
.param tc2_0=1.6539e-07  tc2_w=1.2637e-08
.param jct_0=-0.0460444710839901  jct_w=-1.8e-2 jct_n=4.3569e-05
.param delta_t='temper - 25'
.param lum='l*scale*1e6'   wum='w*scale*1e6'   nsqr='l/w'
.param tc1='tc1_0 + tc1_w * min(wum, 5)'   tc2='tc2_0 + tc2_w * min(wum, 10)'
.param jct='jct_0 + jct_w * min(wum, 2) + jct_n * min(nsqr, 1142.85714285714)'
.param jc1='max(0, (jc1_0 + jc1_w * min(wum, 4) + jc1_n * min(nsqr, 1142.85714285714) + jct * delta_t) / (lum-dl) / (lum-dl))'
.param jc1_r='jc1'
.param tfac='1 + tc1 * delta_t + tc2 * delta_t * delta_t'
.param ro='max(1e-2,rsh/multi*(lum-dl)/(wum-dw))*tfac*(1+factmis)'
rmain n1 n2 'ro*(2-1/(1+jc1_r*v(n1,n2)*v(n1,n2)))'
.ends rppolys
.subckt rnwod n1 n2 l=length w=width  scale='scale_res' multi=1
.param rsh=r_rnwod
.param dw=0.135u
.param pt='temper'
.param pvc1='(1.993e-08/(max(w*scale*1e6, 1.8))+1.259e-09)*(min(l*scale*1e6, 50))+(-5.381e-08/(max(w*scale*1e6, 1.8))+6.448e-08)'   pvc2=0
.param ptc1=1.951e-03   ptc2=8.526e-06
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
.param rmain='rsh/multi*l*scale/(w*scale-dw)*tfac'
.param rend='rend_rnwod'
rn1 n1 1 'rend/multi/(w*scale+0.5u)'
r1 1 2 'max(min(rmain*(1+pvc1*(abs(v(2,1))/l/scale)+pvc2*(v(2,1)/l/scale)*(v(2,1)/l/scale)), rmain*1.5), rmain/2)'
rn2 2 n2 'rend/multi/(w*scale+0.5u)'
.ends rnwod
.subckt rnwsti n1 n2 l=length w=width  scale='scale_res' multi=1
.param rsh=r_rnwsti
.param dw=3.68e-7
.param pt='temper'
.param pvc1='(3.369e-08/(max(w*scale*1e6, 1.8))+8.881e-10)*(min(l*scale*1e6, 50))+(-1.492e-07/(max(w*scale*1e6, 1.8))+1.8e-07)'   pvc2=0
.param ptc1=2.806e-03   ptc2=8.932e-06
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
.param rmain='rsh/multi*l*scale/(w*scale-dw)*tfac'
.param rend='rend_rnwsti'
rn1 n1 1 'rend/multi/(w*scale)'
r1 1 2 'max(min(rmain*(1+pvc1*(abs(v(2,1))/l/scale)+pvc2*(v(2,1)/l/scale)*(v(2,1)/l/scale)), rmain*1.5), rmain/2)'
rn2 2 n2 'rend/multi/(w*scale)'
.ends rnwsti
.subckt rm1l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm1l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6496e-03   ptc2=-5.7895e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm1l
.subckt rm1s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm1s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.3100e-03   ptc2=-5.0480e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm1s
.subckt rm1w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm1w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9890e-03   ptc2=-6.4756e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm1w
.subckt rm2l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm2l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm2l
.subckt rm2s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm2s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm2s
.subckt rm2w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm2w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm2w
.subckt rm3l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm3l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm3l
.subckt rm3s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm3s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm3s
.subckt rm3w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm3w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm3w
.subckt rm4l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm4l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm4l
.subckt rm4s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm4s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm4s
.subckt rm4w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm4w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm4w
.subckt rm5l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm5l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm5l
.subckt rm5s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm5s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm5s
.subckt rm5w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm5w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm5w
.subckt rm6l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm6l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm6l
.subckt rm6s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm6s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm6s
.subckt rm6w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm6w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm6w
.subckt rm7l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm7l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm7l
.subckt rm7s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm7s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm7s
.subckt rm7w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm7w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm7w
.subckt rm8l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm8l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm8l
.subckt rm8s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm8s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm8s
.subckt rm8w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm8w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm8w
.subckt rm9l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm9l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6681e-03   ptc2=-9.5974e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm9l
.subckt rm9s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm9s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6629e-03   ptc2=-9.5672e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm9s
.subckt rm9w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm9w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.8257e-03   ptc2=-1.0493e-06
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm9w
.subckt rm10l n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm10l
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6681e-03   ptc2=-9.5974e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm10l
.subckt rm10s n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm10s
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6629e-03   ptc2=-9.5672e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm10s
.subckt rm10w n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm10w
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.8257e-03   ptc2=-1.0493e-06
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm10w
.subckt rm11 n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rm11
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.8900e-03   ptc2=-1.5000e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rm11
.subckt rmxl n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmxl
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.6617e-03   ptc2=-5.6916e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmxl
.subckt rmxs n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmxs
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.1670e-03   ptc2=-4.7990e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmxs
.subckt rmxw n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmxw
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9415e-03   ptc2=-6.2906e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmxw
.subckt rmyl n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmyl
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.1016e-03   ptc2=-7.4387e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmyl
.subckt rmys n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmys
.param dw=0
.param pvc1=0   pvc2=0   ptc1=2.9413e-03   ptc2=-7.0980e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmys
.subckt rmyw n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmyw
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.4477e-03   ptc2=-9.1619e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmyw
.subckt rmytl n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmytl
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.2086e-03   ptc2=-7.1885e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmytl
.subckt rmyts n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmyts
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.0182e-03   ptc2=-6.4415e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmyts
.subckt rmytw n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmytw
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.5742e-03   ptc2=-8.8010e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmytw
.subckt rmzl n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmzl
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6681e-03   ptc2=-9.5974e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmzl
.subckt rmzs n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmzs
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6629e-03   ptc2=-9.5672e-07
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmzs
.subckt rmzw n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmzw
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.8257e-03   ptc2=-1.0493e-06
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmzw
.subckt rmrl n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmrl
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6620e-03   ptc2=-1.6130e-06
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmrl
.subckt rmrs n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmrs
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6620e-03   ptc2=-1.6130e-06
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmrs
.subckt rmrw n1 n2 l=length w=width scale='scale_res' multi=1
.param rsh=r_rmrw
.param dw=0
.param pvc1=0   pvc2=0   ptc1=3.6620e-03   ptc2=-1.6130e-06
.param pt='temper'
.param tfac='1.0+ptc1*(pt-25.0)+ptc2*(pt-25.0)*(pt-25.0)'
r1 n1 n2 'rsh/multi*l*scale/(w*scale-dw)*(1+pvc1*(abs(v(n2,n1))/l/scale)+pvc2*(v(n2,n1)/l/scale)*(v(n2,n1)/l/scale))*tfac'
.ends rmrw
.param mismatchflag_bip=0
.param mismatchflag_bip_npn=0
.param mismatchflag_disres=0
.param mismatchflag_res=0
.temp "40"
.param sim_temp="40"
.param wireopt=3
.option geoshrink=0.9
.param ccoflag=1
.param ccoflag_12=1
.param ccoflag_18=1
.param ccoflag_18ud15=1
.param ccoflag_cap=1
.param ccoflag_cap_12=1
.param ccoflag_cap_18=1
.param ccoflag_hia=1
.param ccoflag_hvt=1
.param ccoflag_lvt=1
.param ccoflag_na=1
.param ccoflag_na12=1
.param ccoflag_na18=1
.param ccoflag_na18ud15=1
.param rcoflag=1
.param rcoflag_12=1
.param rcoflag_18=1
.param rcoflag_18ud15=1
.param rcoflag_hia=1
.param rcoflag_hvt=1
.param rcoflag_lvt=1
.param rcoflag_na=1
.param rcoflag_na12=1
.param rcoflag_na18=1
.param rcoflag_na18ud15=1
.param rgflag=1
.param rgflag_12=1
.param rgflag_18=1
.param rgflag_18ud15=1
.param rgflag_hia=1
.param rgflag_hvt=1
.param rgflag_lvt=1
.param rgflag_na=1
.param rgflag_na12=1
.param rgflag_na18=1
.param rgflag_na18ud15=1
.subckt od12i VDD VREG emeas_odvref esel_odvref pad rxen rxoutB vrefsel[3] vrefsel[2] vrefsel[1] vrefsel[0] pwrn
.subckt sc_invx2l a y inh_vdd inh_vss
XN0 y a inh_vss inh_vss nch_lvt_mac l=40n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=201.53800n sb=201.53800n sca=2.81171 scb=0.000664299 scc=1.04238e-06 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XP0 y a inh_vdd inh_vdd pch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
.ends sc_invx2l
.subckt cmos12oLS in out outb vddio inh_vdd inh_vss
XM0 outb in inh_vss inh_vss nch_12_mac l=70n w=800n multi=1 nf=1 sd=160.0n ad=1.12e-13 as=1.12e-13 pd=1.88u ps=1.88u nrd=0.029080 nrs=0.029080 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM1 out inb inh_vss inh_vss nch_12_mac l=70n w=800n multi=1 nf=1 sd=160.0n ad=1.12e-13 as=1.12e-13 pd=1.88u ps=1.88u nrd=0.029080 nrs=0.029080 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3 net030 out vddio vddio pch_12_mac l=70n w=2.2u multi=1 nf=2 sd=160.0n ad=1.76e-13 as=3.08e-13 pd=2.52u ps=4.96u nrd=0.014537 nrs=0.014537 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM2 net029 outb vddio vddio pch_12_mac l=70n w=2.2u multi=1 nf=2 sd=160.0n ad=1.76e-13 as=3.08e-13 pd=2.52u ps=4.96u nrd=0.014537 nrs=0.014537 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM5 out inb net029 vddio pch_12_mac l=70n w=2.2u multi=1 nf=2 sd=160.0n ad=1.76e-13 as=3.08e-13 pd=2.52u ps=4.96u nrd=0.014537 nrs=0.014537 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM4 outb in net030 vddio pch_12_mac l=70n w=2.2u multi=1 nf=2 sd=160.0n ad=1.76e-13 as=3.08e-13 pd=2.52u ps=4.96u nrd=0.014537 nrs=0.014537 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XU0 in inb inh_vdd inh_vss sc_invx2l
.ends cmos12oLS
.subckt sc_invx4r a y inh_vdd inh_vss
XP0 y a inh_vdd inh_vdd pch_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.7800n sb=309.7800n sca=10.2911 scb=0.00915362 scc=0.000801174 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=1.47532u enx1=1.46621u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.50641u rey=921.12900n dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=711.5400n
XN0 y a inh_vss inh_vss nch_mac l=40n w=1.32u multi=1 nf=4 sd=160.0n ad=1.056e-13 as=1.452e-13 pd=1.96u ps=2.86u nrd=0.026879 nrs=0.026879 sa=309.7800n sb=309.7800n sca=2.73049 scb=0.000664286 scc=1.04238e-06 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=2.28388u enx1=2.27814u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.28079u rey=1.83014u dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=901.74200n
.ends sc_invx4r
.subckt sc_invx96r a y inh_vdd inh_vss
XN0 y a inh_vss inh_vss nch_mac l=40n w=31.680u multi=1 nf=96 sd=160.0n ad=2.5344e-12 as=2.574e-12 pd=47.040u ps=47.940u nrd=0.001300 nrs=0.001300 sa=3.45041u sb=3.45041u sca=2.31943 scb=0.000664272 scc=1.04238e-06 sa1=632.91500n sa2=1.69248u sa3=1.71443u sa4=3.32594u sb1=632.91500n sb2=1.69248u sb3=1.71443u spa=160.38600n spa1=160.37100n spa2=160.27400n spa3=160.31100n sap=455.79500n spba=181.46200n spba1=183.26500n enx=8.93285u enx1=7.97751u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=8.00925u rey=1.83014u dfm_flag=0 sapb=421.88300n sa5=3.89472u sa6=1.63575u sodx=140.0n sodx1=1.3097u sodx2=2.24258u sody=901.74200n
XP0 y a inh_vdd inh_vdd pch_mac l=40n w=63.360u multi=1 nf=96 sd=160.0n ad=5.0688e-12 as=5.148e-12 pd=78.720u ps=80.280u nrd=0.000966 nrs=0.000966 sa=3.45041u sb=3.45041u sca=9.25666 scb=0.0091425 scc=0.000801174 sa1=632.91500n sa2=1.69248u sa3=1.71443u sa4=3.32594u sb1=632.91500n sb2=1.69248u sb3=1.71443u spa=160.38600n spa1=160.37100n spa2=160.27400n spa3=160.31100n sap=455.79500n spba=181.46200n spba1=183.26500n enx=7.7392u enx1=6.59005u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=9.551u rey=921.12900n dfm_flag=0 sapb=421.88300n sa5=3.89472u sa6=1.63575u sodx=140.0n sodx1=1.3097u sodx2=2.24258u sody=711.5400n
.ends sc_invx96r
.subckt sc_invx20r a y inh_vdd inh_vss
XN0 y a inh_vss inh_vss nch_mac l=40n w=6.6u multi=1 nf=20 sd=160.0n ad=5.28e-13 as=5.676e-13 pd=9.8u ps=10.70u nrd=0.006079 nrs=0.006079 sa=986.10400n sb=986.10400n sca=2.47556 scb=0.000664274 scc=1.04238e-06 sa1=373.62300n sa2=739.82300n sa3=972.17800n sa4=948.90900n sb1=373.62300n sb2=739.82300n sb3=972.17800n spa=161.85700n spa1=161.7900n spa2=161.33500n spa3=161.50600n sap=303.80700n spba=182.85700n spba1=184.66200n enx=3.6282u enx1=3.53155u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=5.32941u rey=1.83014u dfm_flag=0 sapb=313.47300n sa5=1.11825u sa6=932.06900n sodx=140.0n sodx1=595.88400n sodx2=1.43537u sody=901.74200n
XP0 y a inh_vdd inh_vdd pch_mac l=40n w=13.20u multi=1 nf=20 sd=160.0n ad=1.056e-12 as=1.1352e-12 pd=16.40u ps=17.960u nrd=0.004515 nrs=0.004515 sa=986.10400n sb=986.10400n sca=9.57767 scb=0.00914434 scc=0.000801174 sa1=373.62300n sa2=739.82300n sa3=972.17800n sa4=948.90900n sb1=373.62300n sb2=739.82300n sb3=972.17800n spa=161.85700n spa1=161.7900n spa2=161.33500n spa3=161.50600n sap=303.80700n spba=182.85700n spba1=184.66200n enx=2.74175u enx1=2.61013u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=6.01163u rey=921.12900n dfm_flag=0 sapb=313.47300n sa5=1.11825u sa6=932.06900n sodx=140.0n sodx1=595.88400n sodx2=1.43537u sody=711.5400n
.ends sc_invx20r
.subckt cxfr D GN GP S inh_vdd inh_vss nl=40n nw=140n nf=1 pl=40n pw=140n pf=1
XM1 S GN D inh_vss nch_mac l=nl w='nw*nf' multi=1 nf=nf sd=160.0n ad='((nf-int(nf/2)*2)*((140e-9+((nf-1)*160e-9)/2)+0)+((nf+1)-int((nf+1)/2)*2)*((nf/2)*160e-9))*nw' as='((nf-int(nf/2)*2)*((140e-9+((nf-1)*160e-9)/2)+0)+((nf+1)-int((nf+1)/2)*2)*(((280e-9+(nf/2-1)*160e-9)+0)+0))*nw' pd='(nf-int(nf/2)*2)*(((140e-9+((nf-1)*160e-9)/2)+0)*2+(nf+1)*nw)+((nf+1)-int((nf+1)/2)*2)*(((nf/2)*160e-9)*2+nf*nw)' ps='(nf-int(nf/2)*2)*(((140e-9+((nf-1)*160e-9)/2)+0)*2+(nf+1)*nw)+((nf+1)-int((nf+1)/2)*2)*((((280e-9+(nf/2-1)*160e-9)+0)+0)*2+(nf+2)*nw)' sca='((((1e-12/nl)*((0+(1/(2e-6+0*(nl+160e-9))-1/((2e-6+0*(nl+160e-9))+nl)))+(1/(2e-6+0*(nl+160e-9))-1/((2e-6+0*(nl+160e-9))+nl))))/1.0+(1e-12/nw)*(505.050505050505e3-1/(1.98e-6+nw)))+(1e-12/nw)*(1.5625e6-1/(640e-9+nw)))/810e-3' scb='(((0+(1/nl)*(((2e-6+0*(nl+160e-9))/10.0+11.1111e-9)*exp((2e-6+0*(nl+160e-9))*(-9e6))-(((2e-6+0*(nl+160e-9))+nl)/10.0+11.1111e-9)*exp(((2e-6+0*(nl+160e-9))+nl)*(-9e6))))+(1/nl)*(((2e-6+0*(nl+160e-9))/10.0+11.1111e-9)*exp((2e-6+0*(nl+160e-9))*(-9e6))-(((2e-6+0*(nl+160e-9))+nl)/10.0+11.1111e-9)*exp(((2e-6+0*(nl+160e-9))+nl)*(-9e6))))/1.0+(1/nw)*(75.1111e-9*exp(-5.76)-((640e-9+nw)/10.0+11.1111e-9)*exp((640e-9+nw)*(-9e6))))+(1/nw)*(209.1111e-9*exp(-17.82)-((1.98e-6+nw)/10.0+11.1111e-9)*exp((1.98e-6+nw)*(-9e6)))' scc='(((1/nl)*((((0+((2e-6+0*(nl+160e-9))/20.0+2.77778e-9)*exp((2e-6+0*(nl+160e-9))*(-18e6)))-(((2e-6+0*(nl+160e-9))+nl)/20.0+2.77778e-9)*exp(((2e-6+0*(nl+160e-9))+nl)*(-18e6)))+((2e-6+0*(nl+160e-9))/20.0+2.77778e-9)*exp((2e-6+0*(nl+160e-9))*(-18e6)))-(((2e-6+0*(nl+160e-9))+nl)/20.0+2.77778e-9)*exp(((2e-6+0*(nl+160e-9))+nl)*(-18e6))))/1.0+(1/nw)*(34.77778e-9*exp(-11.52)-((640e-9+nw)/20.0+2.77778e-9)*exp((640e-9+nw)*(-18e6))))+(1/nw)*(101.77778e-9*exp(-35.64)-((1.98e-6+nw)/20.0+2.77778e-9)*exp((1.98e-6+nw)*(-18e6)))' dfm_flag=0
XM0 S GP D inh_vdd pch_mac l=pl w='pw*pf' multi=1 nf=pf sd=160.0n ad='((pf-int(pf/2)*2)*((140e-9+((pf-1)*160e-9)/2)+0)+((pf+1)-int((pf+1)/2)*2)*((pf/2)*160e-9))*pw' as='((pf-int(pf/2)*2)*((140e-9+((pf-1)*160e-9)/2)+0)+((pf+1)-int((pf+1)/2)*2)*(((280e-9+(pf/2-1)*160e-9)+0)+0))*pw' pd='(pf-int(pf/2)*2)*(((140e-9+((pf-1)*160e-9)/2)+0)*2+(pf+1)*pw)+((pf+1)-int((pf+1)/2)*2)*(((pf/2)*160e-9)*2+pf*pw)' ps='(pf-int(pf/2)*2)*(((140e-9+((pf-1)*160e-9)/2)+0)*2+(pf+1)*pw)+((pf+1)-int((pf+1)/2)*2)*((((280e-9+(pf/2-1)*160e-9)+0)+0)*2+(pf+2)*pw)' sca='((((1e-12/pl)*((0+(1/(1.2e-6+0*(pl+160e-9))-1/((1.2e-6+0*(pl+160e-9))+pl)))+(1/(1.2e-6+0*(pl+160e-9))-1/((1.2e-6+0*(pl+160e-9))+pl))))/1.0+(1e-12/pw)*(5.88235294117647e6-1/(170e-9+pw)))+(1e-12/pw)*(684.931506849315e3-1/(1.46e-6+pw)))/810e-3' scb='(((0+(1/pl)*(((1.2e-6+0*(pl+160e-9))/10.0+11.1111e-9)*exp((1.2e-6+0*(pl+160e-9))*(-9e6))-(((1.2e-6+0*(pl+160e-9))+pl)/10.0+11.1111e-9)*exp(((1.2e-6+0*(pl+160e-9))+pl)*(-9e6))))+(1/pl)*(((1.2e-6+0*(pl+160e-9))/10.0+11.1111e-9)*exp((1.2e-6+0*(pl+160e-9))*(-9e6))-(((1.2e-6+0*(pl+160e-9))+pl)/10.0+11.1111e-9)*exp(((1.2e-6+0*(pl+160e-9))+pl)*(-9e6))))/1.0+(1/pw)*(157.1111e-9*exp(-13.14)-((1.46e-6+pw)/10.0+11.1111e-9)*exp((1.46e-6+pw)*(-9e6))))+(1/pw)*(28.1111e-9*exp(-1.53)-((170e-9+pw)/10.0+11.1111e-9)*exp((170e-9+pw)*(-9e6)))' scc='(((1/pl)*((((0+((1.2e-6+0*(pl+160e-9))/20.0+2.77778e-9)*exp((1.2e-6+0*(pl+160e-9))*(-18e6)))-(((1.2e-6+0*(pl+160e-9))+pl)/20.0+2.77778e-9)*exp(((1.2e-6+0*(pl+160e-9))+pl)*(-18e6)))+((1.2e-6+0*(pl+160e-9))/20.0+2.77778e-9)*exp((1.2e-6+0*(pl+160e-9))*(-18e6)))-(((1.2e-6+0*(pl+160e-9))+pl)/20.0+2.77778e-9)*exp(((1.2e-6+0*(pl+160e-9))+pl)*(-18e6))))/1.0+(1/pw)*(75.77778e-9*exp(-26.28)-((1.46e-6+pw)/20.0+2.77778e-9)*exp((1.46e-6+pw)*(-18e6))))+(1/pw)*(11.27778e-9*exp(-3.06)-((170e-9+pw)/20.0+2.77778e-9)*exp((170e-9+pw)*(-18e6)))' dfm_flag=0
.ends cxfr
.subckt switch_12_import clk clkb in out pvdd inh_vss
XM0 out clk in inh_vss nch_12_mac l=70n w=2.4u multi=1 nf=4 sd=160.0n ad=1.92e-13 as=2.64e-13 pd=3.04u ps=4.48u nrd=0.012218 nrs=0.012218 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=202.288n spba1=205.319n dfm_flag=0 sapb=244.426n
XM1 out clkb in pvdd pch_12_mac l=70n w=4.8u multi=1 nf=8 sd=160.0n ad=3.84e-13 as=4.56e-13 pd=6.08u ps=7.52u nrd=0.009782 nrs=0.009782 sa=545.317n sb=545.317n sa1=279.161n sa2=472.77n sa3=691.591n sa4=511.925n sb1=279.161n sb2=472.77n sb3=691.591n spa=164.669n spa1=164.513n spa2=163.442n spa3=163.91n sap=251.492n spba=198.962n spba1=201.956n dfm_flag=0 sapb=276.979n
.ends switch_12_import
.subckt sc_invx1_12 a y inh_vdd inh_vss
XM8 y a inh_vss inh_vss nch_12_mac l=70n w=330.0n multi=1 nf=1 sd=160.0n ad=4.62e-14 as=4.62e-14 pd=940.0n ps=940.0n nrd=0.074972 nrs=0.074972 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=886.9n spba1=887.7n dfm_flag=0 sapb=1.668u
XM5 y a inh_vdd inh_vdd pch_12_mac l=70n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.055711 nrs=0.055711 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=886.9n spba1=887.7n dfm_flag=0 sapb=1.668u
.ends sc_invx1_12
.subckt ana_mux_import a b out pvdd sa inh_vss
XI1 selb sela b out pvdd inh_vss switch_12_import
XI0 sela selb a out pvdd inh_vss switch_12_import
XU1 selb sela pvdd inh_vss sc_invx1_12
XU0 sa selb pvdd inh_vss sc_invx1_12
.ends ana_mux_import
.subckt vrefgen_error_in_dec d0 d1 d10 d11 d12 d13 d14 d15 d2 d3 d4 d5 d6 d7 d8 d9 out pvdd s0 s1 s2 s3 inh_vss
XI14 net50 net031 out pvdd s3 inh_vss ana_mux_import
XI13 net44 net43 net031 pvdd s2 inh_vss ana_mux_import
XI12 net46 net45 net50 pvdd s2 inh_vss ana_mux_import
XI11 net32 net31 net43 pvdd s1 inh_vss ana_mux_import
XI10 net34 net33 net44 pvdd s1 inh_vss ana_mux_import
XI9 net36 net35 net45 pvdd s1 inh_vss ana_mux_import
XI8 net38 net37 net46 pvdd s1 inh_vss ana_mux_import
XI7 d7 d6 net34 pvdd s0 inh_vss ana_mux_import
XI6 d3 d2 net32 pvdd s0 inh_vss ana_mux_import
XI5 d1 d0 net31 pvdd s0 inh_vss ana_mux_import
XI4 d5 d4 net33 pvdd s0 inh_vss ana_mux_import
XI3 d11 d10 net36 pvdd s0 inh_vss ana_mux_import
XI2 d9 d8 net35 pvdd s0 inh_vss ana_mux_import
XI1 d13 d12 net37 pvdd s0 inh_vss ana_mux_import
XI0 d15 d14 net38 pvdd s0 inh_vss ana_mux_import
.ends vrefgen_error_in_dec
.subckt sc_invx1r a y inh_vdd inh_vss
XN0 y a inh_vss inh_vss nch_mac l=40n w=330.0n multi=1 nf=1 sd=160.0n ad=4.62e-14 as=4.62e-14 pd=940.0n ps=940.0n nrd=0.074972 nrs=0.074972 sa=140.0n sb=140.0n sca=2.86377 scb=0.000664318 scc=1.04238e-06 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=2u enx1=2u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.0111u rey=1.83014u dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=901.74200n
XP0 y a inh_vdd inh_vdd pch_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.055711 nrs=0.055711 sa=140.0n sb=140.0n sca=10.8078 scb=0.0091796 scc=0.000801174 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=1.2u enx1=1.2u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.07718u rey=921.12900n dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=711.5400n
.ends sc_invx1r
.subckt ls_12 d pvdd q qb vreg inh_vss
XM1 net06 net8 pvdd pvdd pch_12_mac l=70n w=800n multi=1 nf=2 sd=160.0n ad=6.4e-14 as=1.12e-13 pd=1.12u ps=2.16u nrd=0.037591 nrs=0.037591 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM0 net8 net06 pvdd pvdd pch_12_mac l=70n w=800n multi=1 nf=2 sd=160.0n ad=6.4e-14 as=1.12e-13 pd=1.12u ps=2.16u nrd=0.037591 nrs=0.037591 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM3 net06 dbb inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM2 net8 db inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XU1 d db vreg inh_vss sc_invx1r
XU2 db dbb vreg inh_vss sc_invx1r
XU5 net06 q pvdd inh_vss sc_invx1_12
XU3 net8 qb pvdd inh_vss sc_invx1_12
.ends ls_12
.subckt sc_invx4_12 a y inh_vdd inh_vss
XM8 y a inh_vss inh_vss nch_12_mac l=70n w=1.32u multi=1 nf=4 sd=160.0n ad=1.056e-13 as=1.452e-13 pd=1.96u ps=2.86u nrd=0.026879 nrs=0.026879 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=210.3n spba1=213.4n dfm_flag=0 sapb=323n
XM5 y a inh_vdd inh_vdd pch_12_mac l=70n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=210.3n spba1=213.4n dfm_flag=0 sapb=323n
.ends sc_invx4_12
.subckt sc_invx16_12 a y inh_vdd inh_vss
XM8 y a inh_vss inh_vss nch_12_mac l=70n w=5.28u multi=1 nf=16 sd=160.0n ad=4.224e-13 as=4.62e-13 pd=7.84u ps=8.74u nrd=0.007538 nrs=0.007538 sa=921.475n sb=921.475n sa1=353.378n sa2=702.745n sa3=930.644n sa4=860.283n sb1=353.378n sb2=702.745n sb3=930.644n spa=162.323n spa1=162.241n spa2=161.686n spa3=161.926n sap=295.864n spba=199n spba1=201.9n dfm_flag=0 sapb=370.7n
XM5 y a inh_vdd inh_vdd pch_12_mac l=70n w=8.96u multi=1 nf=16 sd=160.0n ad=7.168e-13 as=7.84e-13 pd=11.52u ps=12.88u nrd=0.004750 nrs=0.004750 sa=921.475n sb=921.475n sa1=353.378n sa2=702.745n sa3=930.644n sa4=860.283n sb1=353.378n sb2=702.745n sb3=930.644n spa=162.323n spa1=162.241n spa2=161.686n spa3=161.926n sap=295.864n spba=199n spba1=201.9n dfm_flag=0 sapb=370.7n
.ends sc_invx16_12
.subckt vrefgen_error_in da_0 da_1 da_2 da_3 out powerdown pvdd vreg inh_vss
XXR2 a15 a14 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR3 a14 a13 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR4 a13 a12 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR5 a12 a11 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR6 a11 a10 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR7 a10 a9 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR8 a9 a8 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR9 a8 a7 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR10 a4 a3 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR11 a5 a4 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR12 a6 a5 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR13 a7 a6 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR14 a3 a2 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR15 a2 a1 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR16 a1 a0 inh_vss rppolywo_m lr=1u wr=1u multi=1 m=1
XXR1_1__dmy0 net019 XR1_1__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_2__dmy0 XR1_1__dmy0 XR1_2__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_3__dmy0 XR1_2__dmy0 XR1_3__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_4__dmy0 XR1_3__dmy0 XR1_4__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_5__dmy0 XR1_4__dmy0 XR1_5__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_6__dmy0 XR1_5__dmy0 XR1_6__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_7__dmy0 XR1_6__dmy0 XR1_7__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_8__dmy0 XR1_7__dmy0 XR1_8__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_9__dmy0 XR1_8__dmy0 XR1_9__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_10__dmy0 XR1_9__dmy0 XR1_10__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_11__dmy0 XR1_10__dmy0 XR1_11__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_12__dmy0 XR1_11__dmy0 XR1_12__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_13__dmy0 XR1_12__dmy0 XR1_13__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_14__dmy0 XR1_13__dmy0 XR1_14__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_15__dmy0 XR1_14__dmy0 XR1_15__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_16__dmy0 XR1_15__dmy0 XR1_16__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_17__dmy0 XR1_16__dmy0 XR1_17__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_18__dmy0 XR1_17__dmy0 XR1_18__dmy0 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR1_19__dmy0 XR1_18__dmy0 a15 inh_vss rppolywo_m lr=1.04u wr=1u multi=1 m=1
XXR0_1__dmy0 a0 XR0_1__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_2__dmy0 XR0_1__dmy0 XR0_2__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_3__dmy0 XR0_2__dmy0 XR0_3__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_4__dmy0 XR0_3__dmy0 XR0_4__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_5__dmy0 XR0_4__dmy0 XR0_5__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_6__dmy0 XR0_5__dmy0 XR0_6__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_7__dmy0 XR0_6__dmy0 XR0_7__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_8__dmy0 XR0_7__dmy0 XR0_8__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_9__dmy0 XR0_8__dmy0 XR0_9__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_10__dmy0 XR0_9__dmy0 XR0_10__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_11__dmy0 XR0_10__dmy0 XR0_11__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_12__dmy0 XR0_11__dmy0 XR0_12__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_13__dmy0 XR0_12__dmy0 XR0_13__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_14__dmy0 XR0_13__dmy0 XR0_14__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_15__dmy0 XR0_14__dmy0 XR0_15__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_16__dmy0 XR0_15__dmy0 XR0_16__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_17__dmy0 XR0_16__dmy0 XR0_17__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_18__dmy0 XR0_17__dmy0 XR0_18__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_19__dmy0 XR0_18__dmy0 XR0_19__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_20__dmy0 XR0_19__dmy0 XR0_20__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_21__dmy0 XR0_20__dmy0 XR0_21__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_22__dmy0 XR0_21__dmy0 XR0_22__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_23__dmy0 XR0_22__dmy0 XR0_23__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_24__dmy0 XR0_23__dmy0 XR0_24__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_25__dmy0 XR0_24__dmy0 XR0_25__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_26__dmy0 XR0_25__dmy0 XR0_26__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_27__dmy0 XR0_26__dmy0 XR0_27__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_28__dmy0 XR0_27__dmy0 XR0_28__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_29__dmy0 XR0_28__dmy0 XR0_29__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_30__dmy0 XR0_29__dmy0 XR0_30__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_31__dmy0 XR0_30__dmy0 XR0_31__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_32__dmy0 XR0_31__dmy0 XR0_32__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_33__dmy0 XR0_32__dmy0 XR0_33__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_34__dmy0 XR0_33__dmy0 XR0_34__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_35__dmy0 XR0_34__dmy0 XR0_35__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_36__dmy0 XR0_35__dmy0 XR0_36__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_37__dmy0 XR0_36__dmy0 XR0_37__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_38__dmy0 XR0_37__dmy0 XR0_38__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_39__dmy0 XR0_38__dmy0 XR0_39__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_40__dmy0 XR0_39__dmy0 XR0_40__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_41__dmy0 XR0_40__dmy0 XR0_41__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_42__dmy0 XR0_41__dmy0 XR0_42__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_43__dmy0 XR0_42__dmy0 XR0_43__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_44__dmy0 XR0_43__dmy0 XR0_44__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_45__dmy0 XR0_44__dmy0 XR0_45__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_46__dmy0 XR0_45__dmy0 XR0_46__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_47__dmy0 XR0_46__dmy0 XR0_47__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_48__dmy0 XR0_47__dmy0 XR0_48__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_49__dmy0 XR0_48__dmy0 XR0_49__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_50__dmy0 XR0_49__dmy0 XR0_50__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_51__dmy0 XR0_50__dmy0 XR0_51__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_52__dmy0 XR0_51__dmy0 XR0_52__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_53__dmy0 XR0_52__dmy0 XR0_53__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_54__dmy0 XR0_53__dmy0 XR0_54__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_55__dmy0 XR0_54__dmy0 XR0_55__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_56__dmy0 XR0_55__dmy0 XR0_56__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_57__dmy0 XR0_56__dmy0 XR0_57__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_58__dmy0 XR0_57__dmy0 XR0_58__dmy0 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XXR0_59__dmy0 XR0_58__dmy0 net024 inh_vss rppolywo_m lr=1.005u wr=1u multi=1 m=1
XI4 a0 a1 a10 a11 a12 a13 a14 a15 a2 a3 a4 a5 a6 a7 a8 a9 out pvdd s0 s1 s2 s3 inh_vss vrefgen_error_in_dec
XI6 da_2 pvdd net09 net014 vreg inh_vss ls_12
XI5 da_3 pvdd net012 net013 vreg inh_vss ls_12
XI7 da_1 pvdd net07 net08 vreg inh_vss ls_12
XI16 powerdown pvdd net025 net021 vreg inh_vss ls_12
XI8 da_0 pvdd net04 net03 vreg inh_vss ls_12
XU0 net012 net011 pvdd inh_vss sc_invx1_12
XU5 net07 net06 pvdd inh_vss sc_invx1_12
XU2 net09 net010 pvdd inh_vss sc_invx1_12
XU6 net04 net05 pvdd inh_vss sc_invx1_12
XM0 net019 pwrdn pvdd pvdd pch_12_mac l=70n w=30u multi=1 nf=30 sd=160.0n ad=2.4e-12 as=2.52e-12 pd=34.8u ps=37.04u nrd=0.001506 nrs=0.001506 sa=1.50916u sb=1.50916u sa1=437.336n sa2=991.492n sa3=1.18243u sa4=1.40782u sb1=437.336n sb2=991.492n sb3=1.18243u spa=161.236n spa1=161.191n spa2=160.891n spa3=161.02n sap=346.278n spba=196.748n spba1=199.717n dfm_flag=0 sapb=358.265n
XM1 net024 pwrdnb inh_vss inh_vss nch_12_mac l=70n w=20u multi=1 nf=20 sd=160.0n ad=1.6e-12 as=1.72e-12 pd=23.2u ps=25.44u nrd=0.001504 nrs=0.001504 sa=1.09596u sb=1.09596u sa1=381.185n sa2=795.251n sa3=1.01548u sa4=1.02252u sb1=381.185n sb2=795.251n sb3=1.01548u spa=161.857n spa1=161.79n spa2=161.343n spa3=161.536n sap=312.569n spba=197.138n spba1=200.112n dfm_flag=0 sapb=330.374n
XU1 net011 s3 pvdd inh_vss sc_invx4_12
XU4 net06 s1 pvdd inh_vss sc_invx4_12
XU3 net010 s2 pvdd inh_vss sc_invx4_12
XU7 net05 s0 pvdd inh_vss sc_invx4_12
XU8 net025 net028 pvdd inh_vss sc_invx4_12
XU11 net021 net030 pvdd inh_vss sc_invx4_12
XU9 net028 pwrdn pvdd inh_vss sc_invx16_12
XU10 net030 pwrdnb pvdd inh_vss sc_invx16_12
.ends vrefgen_error_in
.subckt eEsdndio pad inh_vss
D0 inh_vss pad ndio_12 area=6e-11 pj=8.3e-05 m=1
.ends eEsdndio
.subckt eEsdpdio pad vtt
D1 pad vtt pdio_12 area=6e-11 pj=8.3e-05 m=1
.ends eEsdpdio
.subckt eEsdhbm pad vtt inh_vss
XI9 pad inh_vss eEsdndio
XI8 pad vtt eEsdpdio
.ends eEsdhbm
.subckt eEsdcdm in out vtt inh_vss
D0 inh_vss out ndio_12 area=4.352e-12 pj=9.12e-06 m=1
XXR0 in out vtt rppolywo_m lr=2u wr=2u multi=5 m=1
D1 out vtt pdio_12 area=4.352e-12 pj=9.12e-06 m=1
.ends eEsdcdm
.subckt sc_invx6_12 a y inh_vdd inh_vss
XM8 y a inh_vss inh_vss nch_12_mac l=70n w=1.98u multi=1 nf=6 sd=160.0n ad=1.584e-13 as=1.98e-13 pd=2.94u ps=3.84u nrd=0.018827 nrs=0.018827 sa=441.862n sb=441.862n sa1=253.113n sa2=398.819n sa3=600.454n sa4=416.572n sb1=253.113n sb2=398.819n sb3=600.454n spa=166.245n spa1=166.045n spa2=164.654n spa3=165.267n sap=236.148n spba=204.723n spba1=207.754n dfm_flag=0 sapb=329.879n
XM5 y a inh_vdd inh_vdd pch_12_mac l=70n w=3.96u multi=1 nf=6 sd=160.0n ad=3.168e-13 as=3.96e-13 pd=4.92u ps=6.48u nrd=0.013983 nrs=0.013983 sa=441.862n sb=441.862n sa1=253.113n sa2=398.819n sa3=600.454n sa4=416.572n sb1=253.113n sb2=398.819n sb3=600.454n spa=166.245n spa1=166.045n spa2=164.654n spa3=165.267n sap=236.148n spba=204.723n spba1=207.754n dfm_flag=0 sapb=329.879n
.ends sc_invx6_12
.subckt sc_invx8r a y inh_vdd inh_vss
XP0 y a inh_vdd inh_vdd pch_mac l=40n w=5.28u multi=1 nf=8 sd=160.0n ad=4.224e-13 as=5.016e-13 pd=6.56u ps=8.12u nrd=0.010760 nrs=0.010760 sa=499.16600n sb=499.16600n sca=9.95574 scb=0.00914783 scc=0.000801174 sa1=274.42700n sa2=442.39700n sa3=656.64400n sa4=482.30100n sb1=274.42700n sb2=442.39700n sb3=656.64400n spa=164.66900n spa1=164.51300n spa2=163.42100n spa3=163.83800n sap=245.63900n spba=185.72100n spba1=187.52900n enx=1.81526u enx1=1.7842u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.97078u rey=921.12900n dfm_flag=0 sapb=269.45200n sa5=558.0500n sa6=634.76800n sodx=140.0n sodx1=397.24900n sodx2=1.11642u sody=711.5400n
XN0 y a inh_vss inh_vss nch_mac l=40n w=2.64u multi=1 nf=8 sd=160.0n ad=2.112e-13 as=2.508e-13 pd=3.92u ps=4.82u nrd=0.014487 nrs=0.014487 sa=499.16600n sb=499.16600n sca=2.62336 scb=0.000664279 scc=1.04238e-06 sa1=274.42700n sa2=442.39700n sa3=656.64400n sa4=482.30100n sb1=274.42700n sb2=442.39700n sb3=656.64400n spa=164.66900n spa1=164.51300n spa2=163.42100n spa3=163.83800n sap=245.63900n spba=185.72100n spba1=187.52900n enx=2.64131u enx1=2.62048u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.59103u rey=1.83014u dfm_flag=0 sapb=269.45200n sa5=558.0500n sa6=634.76800n sodx=140.0n sodx1=397.24900n sodx2=1.11642u sody=901.74200n
.ends sc_invx8r
.subckt sc_nand2x4r a b y inh_vdd inh_vss
XNb net21 b inh_vss inh_vss nch_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.013439 nrs=0.013439 sa=309.7800n sb=309.7800n sca=2.19193 scb=0.000356858 scc=5.23214e-07 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=2.28388u enx1=2.27814u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.28079u rey=1.83014u dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=901.74200n
XNa y a net21 inh_vss nch_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.013439 nrs=0.013439 sa=309.7800n sb=309.7800n sca=2.19193 scb=0.000356858 scc=5.23214e-07 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=2.28388u enx1=2.27814u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.28079u rey=1.83014u dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=901.74200n
XPa y a inh_vdd inh_vdd pch_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.7800n sb=309.7800n sca=10.2911 scb=0.00915362 scc=0.000801174 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=1.47532u enx1=1.46621u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.50641u rey=921.12900n dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=711.5400n
XPb y b inh_vdd inh_vdd pch_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.7800n sb=309.7800n sca=10.2911 scb=0.00915362 scc=0.000801174 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=1.47532u enx1=1.46621u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.50641u rey=921.12900n dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=711.5400n
.ends sc_nand2x4r
.subckt DamNcap1p8x1p8V12 minus plus
XC0 plus minus nmoscap_12 lr=1.8u wr=1.8u multi=1
.ends DamNcap1p8x1p8V12
.subckt cxfr_mv D GN GP S inh_vdd inh_vss nl=70n nw=140n nf=1 nsd=140n pl=70n pw=140n pf=1 psd=140n
XM0 S GN D inh_vss nch_12_mac l=nl w='nw*nf' multi=1 nf=nf sd=nsd ad='((nf-int(nf/2)*2)*((140e-9+((nf-1)*160e-9)/2)+0)+((nf+1)-int((nf+1)/2)*2)*((nf/2)*160e-9))*nw' as='((nf-int(nf/2)*2)*((140e-9+((nf-1)*160e-9)/2)+0)+((nf+1)-int((nf+1)/2)*2)*(((280e-9+(nf/2-1)*160e-9)+0)+0))*nw' pd='(nf-int(nf/2)*2)*(((140e-9+((nf-1)*160e-9)/2)+0)*2+(nf+1)*nw)+((nf+1)-int((nf+1)/2)*2)*(((nf/2)*160e-9)*2+nf*nw)' ps='(nf-int(nf/2)*2)*(((140e-9+((nf-1)*160e-9)/2)+0)*2+(nf+1)*nw)+((nf+1)-int((nf+1)/2)*2)*((((280e-9+(nf/2-1)*160e-9)+0)+0)*2+(nf+2)*nw)' dfm_flag=0
XM1 S GP D inh_vdd pch_12_mac l=pl w='pw*pf' multi=1 nf=pf sd=psd ad='((pf-int(pf/2)*2)*((140e-9+((pf-1)*160e-9)/2)+0)+((pf+1)-int((pf+1)/2)*2)*((pf/2)*160e-9))*pw' as='((pf-int(pf/2)*2)*((140e-9+((pf-1)*160e-9)/2)+0)+((pf+1)-int((pf+1)/2)*2)*(((280e-9+(pf/2-1)*160e-9)+0)+0))*pw' pd='(pf-int(pf/2)*2)*(((140e-9+((pf-1)*160e-9)/2)+0)*2+(pf+1)*pw)+((pf+1)-int((pf+1)/2)*2)*(((pf/2)*160e-9)*2+pf*pw)' ps='(pf-int(pf/2)*2)*(((140e-9+((pf-1)*160e-9)/2)+0)*2+(pf+1)*pw)+((pf+1)-int((pf+1)/2)*2)*((((280e-9+(pf/2-1)*160e-9)+0)+0)*2+(pf+2)*pw)' dfm_flag=0
.ends cxfr_mv
.subckt sc_invx8_12 a y inh_vdd inh_vss
XM8 y a inh_vss inh_vss nch_12_mac l=70n w=2.64u multi=1 nf=8 sd=160n ad=211.2f as=250.8f pd=3.92u ps=4.82u nrd=0.01449 nrs=0.01449 sa=545.3n sb=545.3n sa1=279.2n sa2=472.8n sa3=691.6n sa4=511.9n sb1=279.2n sb2=472.8n sb3=691.6n spa=164.7n spa1=164.5n spa2=163.4n spa3=163.9n sap=251.5n spba=202.3n spba1=205.3n dfm_flag=0 sapb=338.9n
XM5 y a inh_vdd inh_vdd pch_12_mac l=70n w=5.28u multi=1 nf=8 sd=160n ad=422.4f as=501.6f pd=6.56u ps=8.12u nrd=0.01076 nrs=0.01076 sa=545.3n sb=545.3n sa1=279.2n sa2=472.8n sa3=691.6n sa4=511.9n sb1=279.2n sb2=472.8n sb3=691.6n spa=164.7n spa1=164.5n spa2=163.4n spa3=163.9n sap=251.5n spba=202.3n spba1=205.3n dfm_flag=0 sapb=338.9n
.ends sc_invx8_12
.subckt DamNcap2x2p4V12 minus plus
XC1 plus minus nmoscap_12 lr=2u wr=2.4u multi=1
.ends DamNcap2x2p4V12
.subckt sc_invx2_12 a y inh_vdd inh_vss
XM8 y a inh_vss inh_vss nch_12_mac l=70n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=238.3n spba1=241.4n dfm_flag=0 sapb=348.7n
XM5 y a inh_vdd inh_vdd pch_12_mac l=70n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=238.3n spba1=241.4n dfm_flag=0 sapb=348.7n
.ends sc_invx2_12
.subckt cmos12iBias rxen vbiasn vbiasp vdd inh_vdd inh_vss
XM112 vdd vdd vdd vdd pch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM111 vdd vdd vdd vdd pch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM103 vbiasp vbiasp vdd vdd pch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM10 vdd vbiasp vdd vdd pch_12_mac l=900n w=3.6u multi=1 nf=4 sd=160.0n ad=2.88e-13 as=3.96e-13 pd=4.24u ps=6.28u nrd=0.012100 nrs=0.012100 sa=912.755n sb=912.755n sa1=274.265n sa2=676.078n sa3=702.449n sa4=460.647n sb1=274.265n sb2=676.078n sb3=702.449n spa=162.463n spa1=162.444n spa2=162.356n spa3=162.455n sap=236.406n spba=299.854n spba1=353.929n dfm_flag=0 sapb=279.35n
XM108 net0119 rxenb12 vdd vdd pch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM110 vdd vdd vdd vdd pch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM109 vdd vdd vdd vdd pch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM9 vdd net017 vdd vdd pch_12_mac l=1u w=6.3u multi=1 nf=7 sd=160.0n ad=5.58e-13 as=5.58e-13 pd=8.44u ps=8.44u nrd=0.007371 nrs=0.007371 sa=1.70482u sb=1.70482u sa1=358.136n sa2=1.10161u sa3=909.373n sa4=771.86n sb1=358.136n sb2=1.10161u sb3=909.373n spa=161.404n spa1=161.392n spa2=161.339n spa3=161.401n sap=280.284n spba=334.59n spba1=399.555n dfm_flag=0 sapb=321.304n
XM104 vbiasp rxenbb12 vdd vdd pch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM116 inh_vss inh_vss inh_vss inh_vss nch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM115 inh_vss inh_vss inh_vss inh_vss nch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM114 inh_vss inh_vss inh_vss inh_vss nch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM113 inh_vss inh_vss inh_vss inh_vss nch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM105 vbiasn vbiasn inh_vss inh_vss nch_12_mac l=200n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=242.857n sb=242.857n sa1=179.667n sa2=233.669n sa3=356.204n sa4=219.1n sb1=179.667n sb2=233.669n sb3=356.204n spa=164.95n spa1=164.925n spa2=164.73n spa3=164.859n sap=184.41n spba=221.192n spba1=230.208n dfm_flag=0 sapb=231.646n
XM106 net092 rxenbb12 inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM107 vbiasn rxenb12 inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XC0 inh_vss vbiasn DamNcap1p8x1p8V12
XXR5_1__dmy0 net0119 XR5_1__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_2__dmy0 XR5_1__dmy0 XR5_2__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_3__dmy0 XR5_2__dmy0 XR5_3__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_4__dmy0 XR5_3__dmy0 XR5_4__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_5__dmy0 XR5_4__dmy0 XR5_5__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_6__dmy0 XR5_5__dmy0 XR5_6__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_7__dmy0 XR5_6__dmy0 XR5_7__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_8__dmy0 XR5_7__dmy0 XR5_8__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_9__dmy0 XR5_8__dmy0 XR5_9__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_10__dmy0 XR5_9__dmy0 XR5_10__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_11__dmy0 XR5_10__dmy0 XR5_11__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_12__dmy0 XR5_11__dmy0 XR5_12__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_13__dmy0 XR5_12__dmy0 XR5_13__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_14__dmy0 XR5_13__dmy0 XR5_14__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_15__dmy0 XR5_14__dmy0 XR5_15__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_16__dmy0 XR5_15__dmy0 XR5_16__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_17__dmy0 XR5_16__dmy0 XR5_17__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_18__dmy0 XR5_17__dmy0 XR5_18__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_19__dmy0 XR5_18__dmy0 XR5_19__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_20__dmy0 XR5_19__dmy0 vbiasn inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_1__dmy0 vbiasp XR4_1__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_2__dmy0 XR4_1__dmy0 XR4_2__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_3__dmy0 XR4_2__dmy0 XR4_3__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_4__dmy0 XR4_3__dmy0 XR4_4__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_5__dmy0 XR4_4__dmy0 XR4_5__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_6__dmy0 XR4_5__dmy0 XR4_6__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_7__dmy0 XR4_6__dmy0 XR4_7__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_8__dmy0 XR4_7__dmy0 XR4_8__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_9__dmy0 XR4_8__dmy0 XR4_9__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_10__dmy0 XR4_9__dmy0 XR4_10__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_11__dmy0 XR4_10__dmy0 XR4_11__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_12__dmy0 XR4_11__dmy0 XR4_12__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_13__dmy0 XR4_12__dmy0 XR4_13__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_14__dmy0 XR4_13__dmy0 XR4_14__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_15__dmy0 XR4_14__dmy0 XR4_15__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_16__dmy0 XR4_15__dmy0 XR4_16__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_17__dmy0 XR4_16__dmy0 XR4_17__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_18__dmy0 XR4_17__dmy0 XR4_18__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_19__dmy0 XR4_18__dmy0 XR4_19__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_20__dmy0 XR4_19__dmy0 net092 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XU10 inh_vss rxenb12 rxenbb12 net017 vdd inh_vss cxfr_mv m=1 nl=70n nw=1u nf=8 nsd=140.0n pl=70n pw=1u pf=8 psd=140.0n
XU9 vbiasp rxenbb12 rxenb12 net017 vdd inh_vss cxfr_mv m=1 nl=70n nw=1u nf=8 nsd=140.0n pl=70n pw=1u pf=8 psd=140.0n
XU7 vdd rxenb12 rxenbb12 net050 vdd inh_vss cxfr_mv m=1 nl=70n nw=1u nf=8 nsd=140.0n pl=70n pw=1u pf=8 psd=140.0n
XU8 vbiasn rxenbb12 rxenb12 net050 vdd inh_vss cxfr_mv m=1 nl=70n nw=1u nf=8 nsd=140.0n pl=70n pw=1u pf=8 psd=140.0n
XU18 net058 rxenbb12 vdd inh_vss sc_invx8_12
XU19 net0108 rxenb12 vdd inh_vss sc_invx8_12
XU17 net0101 net0108 vdd inh_vss sc_invx8_12
XU0 net0102 net058 vdd inh_vss sc_invx8_12
XC1 inh_vss net050 DamNcap2x2p4V12
XI22_4_ rxen net0102 net0101 vdd inh_vdd inh_vss cmos12oLS
XI22_3_ rxen net0102 net0101 vdd inh_vdd inh_vss cmos12oLS
XI22_2_ rxen net0102 net0101 vdd inh_vdd inh_vss cmos12oLS
XI22_1_ rxen net0102 net0101 vdd inh_vdd inh_vss cmos12oLS
XI22_0_ rxen net0102 net0101 vdd inh_vdd inh_vss cmos12oLS
XU20 net0108 net058 vdd inh_vss sc_invx2_12
XU1 net058 net0108 vdd inh_vss sc_invx2_12
.ends cmos12iBias
.subckt sc_nand2x1r a b y inh_vdd inh_vss
XPa y a inh_vdd inh_vdd pch_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.055711 nrs=0.055711 sa=140.0n sb=140.0n sca=10.8078 scb=0.0091796 scc=0.000801174 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=1.2u enx1=1.2u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.07718u rey=921.12900n dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=711.5400n
XPb y b inh_vdd inh_vdd pch_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.055711 nrs=0.055711 sa=140.0n sb=140.0n sca=10.8078 scb=0.0091796 scc=0.000801174 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=1.2u enx1=1.2u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.07718u rey=921.12900n dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=711.5400n
Xnb net21 b inh_vss inh_vss nch_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.037486 nrs=0.037486 sa=140.0n sb=140.0n sca=2.32522 scb=0.00035689 scc=5.23214e-07 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=2u enx1=2u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.0111u rey=1.83014u dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=901.74200n
XNa y a net21 inh_vss nch_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.037486 nrs=0.037486 sa=140.0n sb=140.0n sca=2.32522 scb=0.00035689 scc=5.23214e-07 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=2u enx1=2u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.0111u rey=1.83014u dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=901.74200n
.ends sc_nand2x1r
.subckt ckRxOffsetN bottom off[3] off[2] off[1] off[0] tiehi top inh_vss
XM3_7_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_6_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_5_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_4_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_3_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_2_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_1_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM3_0_ top off[3] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM2_3_ top off[2] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM2_2_ top off[2] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM2_1_ top off[2] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM2_0_ top off[2] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM1_1_ top off[1] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM1_0_ top off[1] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
Xn5 top tiehi bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
XM0 top off[0] bottom inh_vss nch_12_mac l=70n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=208.495n spba1=211.941n dfm_flag=0 sapb=190.886n
.ends ckRxOffsetN
.subckt ckRxOffsetP bottom off[3] off[2] off[1] off[0] tielo top inh_vdd
XM1_1_ bottom off[1] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM1_0_ bottom off[1] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_7_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_6_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_5_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_4_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_3_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_2_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_1_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM3_0_ bottom off[3] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM2_3_ bottom off[2] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM2_2_ bottom off[2] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM2_1_ bottom off[2] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM2_0_ bottom off[2] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
Xp5 bottom tielo top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM0 bottom off[0] top inh_vdd pch_12_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
.ends ckRxOffsetP
.subckt cmos12iAmpCore VDD in inb offcalen offcalenb offcalenbb offset[4] offset[3] offset[2] offset[1] offset[0] on op pd_rxen rxen inh_vdd inh_vss
XU2 oceniob offcalenbb VDD inh_vss sc_invx6_12
XU1 ocenio offcalenb VDD inh_vss sc_invx6_12
XI7_3_ offp[3] offp12b[3] offp12[3] VDD inh_vdd inh_vss cmos12oLS
XI7_2_ offp[2] offp12b[2] offp12[2] VDD inh_vdd inh_vss cmos12oLS
XI7_1_ offp[1] offp12b[1] offp12[1] VDD inh_vdd inh_vss cmos12oLS
XI7_0_ offp[0] offp12b[0] offp12[0] VDD inh_vdd inh_vss cmos12oLS
XI1_1_ enb eniob enio VDD inh_vdd inh_vss cmos12oLS
XI1_0_ enb eniob enio VDD inh_vdd inh_vss cmos12oLS
XI5_3_ net0141[0] offn12[3] offn12b[3] VDD inh_vdd inh_vss cmos12oLS
XI5_2_ net0141[1] offn12[2] offn12b[2] VDD inh_vdd inh_vss cmos12oLS
XI5_1_ net0141[2] offn12[1] offn12b[1] VDD inh_vdd inh_vss cmos12oLS
XI5_0_ net0141[3] offn12[0] offn12b[0] VDD inh_vdd inh_vss cmos12oLS
Xlsocen_3_ offcalen ocenio oceniob VDD inh_vdd inh_vss cmos12oLS
Xlsocen_2_ offcalen ocenio oceniob VDD inh_vdd inh_vss cmos12oLS
Xlsocen_1_ offcalen ocenio oceniob VDD inh_vdd inh_vss cmos12oLS
Xlsocen_0_ offcalen ocenio oceniob VDD inh_vdd inh_vss cmos12oLS
XU8 enb en inh_vdd inh_vss sc_invx8r
XU7 rxen pd_rxen enb inh_vdd inh_vss sc_nand2x4r
XI16 en vbiasn vbiasp VDD inh_vdd inh_vss cmos12iBias
XU16 offset[4] net283 inh_vdd inh_vss sc_invx1r
XU4_3_ net324[0] net0141[0] inh_vdd inh_vss sc_invx1r
XU4_2_ net324[1] net0141[1] inh_vdd inh_vss sc_invx1r
XU4_1_ net324[2] net0141[2] inh_vdd inh_vss sc_invx1r
XU4_0_ net324[3] net0141[3] inh_vdd inh_vss sc_invx1r
XU3_3_ en net325[0] offp[3] inh_vdd inh_vss sc_nand2x1r
XU3_2_ en net325[1] offp[2] inh_vdd inh_vss sc_nand2x1r
XU3_1_ en net325[2] offp[1] inh_vdd inh_vss sc_nand2x1r
XU3_0_ en net325[3] offp[0] inh_vdd inh_vss sc_nand2x1r
XU12_3_ offset[3] net283 net325[0] inh_vdd inh_vss sc_nand2x1r
XU12_2_ offset[2] net283 net325[1] inh_vdd inh_vss sc_nand2x1r
XU12_1_ offset[1] net283 net325[2] inh_vdd inh_vss sc_nand2x1r
XU12_0_ offset[0] net283 net325[3] inh_vdd inh_vss sc_nand2x1r
XU13_3_ en net323[0] net324[0] inh_vdd inh_vss sc_nand2x1r
XU13_2_ en net323[1] net324[1] inh_vdd inh_vss sc_nand2x1r
XU13_1_ en net323[2] net324[2] inh_vdd inh_vss sc_nand2x1r
XU13_0_ en net323[3] net324[3] inh_vdd inh_vss sc_nand2x1r
XU14_3_ offset[4] offset[3] net323[0] inh_vdd inh_vss sc_nand2x1r
XU14_2_ offset[4] offset[2] net323[1] inh_vdd inh_vss sc_nand2x1r
XU14_1_ offset[4] offset[1] net323[2] inh_vdd inh_vss sc_nand2x1r
XU14_0_ offset[4] offset[0] net323[3] inh_vdd inh_vss sc_nand2x1r
XM36 in offcalenbb inb inh_vss nch_12_mac l=70n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.006649 nrs=0.006649 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=202.288n spba1=205.319n dfm_flag=0 sapb=244.426n
Xinn headin in net075 inh_vss nch_12_mac l=150.0n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.006649 nrs=0.006649 sa=388.666n sb=388.666n sa1=227.236n sa2=354.562n sa3=541.173n sa4=345.184n sb1=227.236n sb2=354.562n sb3=541.173n spa=162.463n spa1=162.444n spa2=162.298n spa3=162.385n sap=212.983n spba=222.403n spba1=228.634n dfm_flag=0 sapb=266.153n
XM3 headref inb net084 inh_vss nch_12_mac l=150.0n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.006649 nrs=0.006649 sa=388.666n sb=388.666n sa1=227.236n sa2=354.562n sa3=541.173n sa4=345.184n sb1=227.236n sb2=354.562n sb3=541.173n spa=162.463n spa1=162.444n spa2=162.298n spa3=162.385n sap=212.983n spba=222.403n spba1=228.634n dfm_flag=0 sapb=266.153n
XM9 headin eniob inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM20 tailn eniob inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM1 net327 enio inh_vss inh_vss nch_12_mac l=70n w=12.0u multi=1 nf=12 sd=160.0n ad=9.6e-13 as=1.08e-12 pd=13.92u ps=16.16u nrd=0.002453 nrs=0.002453 sa=739.143n sb=739.143n sa1=320.464n sa2=597.542n sa3=827.446n sa4=691.15n sb1=320.464n sb2=597.542n sb3=827.446n spa=163.103n spa1=162.995n spa2=162.263n spa3=162.581n sap=276.12n spba=197.934n spba1=200.917n dfm_flag=0 sapb=299.055n
XM0 tailn vbiasn net327 inh_vss nch_12_mac l=200n w=16.0u multi=1 nf=16 sd=160.0n ad=1.28e-12 as=1.4e-12 pd=18.56u ps=20.8u nrd=0.001865 nrs=0.001865 sa=1.30442u sb=1.30442u sa1=377.952n sa2=893.294n sa3=1.06016u sa4=1.06817u sb1=377.952n sb2=893.294n sb3=1.06016u spa=160.613n spa1=160.608n spa2=160.565n spa3=160.593n sap=308.397n spba=248.146n spba1=255.744n dfm_flag=0 sapb=373.804n
XM8 headref eniob inh_vss inh_vss nch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.011617 nrs=0.011617 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XXR2_1__dmy0 op XR2_1__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR2_2__dmy0 XR2_1__dmy0 XR2_2__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR2_3__dmy0 XR2_2__dmy0 inh_vss inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR0_1__dmy0 on XR0_1__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR0_2__dmy0 XR0_1__dmy0 XR0_2__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR0_3__dmy0 XR0_2__dmy0 inh_vss inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
Xoffninb tailn offn12[3] offn12[2] offn12[1] offn12[0] enio net084 inh_vss ckRxOffsetN
Xoffnin tailn offp12[3] offp12[2] offp12[1] offp12[0] enio net075 inh_vss ckRxOffsetN
XM40 in offcalenb inb VDD pch_12_mac l=80n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.009877 nrs=0.009877 sa=338.689n sb=338.689n sa1=221.443n sa2=317.974n sa3=486.769n sa4=319.355n sb1=221.443n sb2=317.974n sb3=486.769n spa=162.463n spa1=162.444n spa2=162.291n spa3=162.366n sap=207.166n spba=200.998n spba1=204.373n dfm_flag=0 sapb=250.308n
XM25 net068 eniob VDD VDD pch_12_mac l=70n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.009877 nrs=0.009877 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=202.288n spba1=205.319n dfm_flag=0 sapb=244.426n
XM11 tailp enio VDD VDD pch_12_mac l=70n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=209.397n sb=209.397n sa1=174.687n sa2=205.977n sa3=286.184n sa4=203.362n sb1=174.687n sb2=205.977n sb3=286.184n spa=179.221n spa1=178.832n spa2=175.794n spa3=177.223n sap=192.81n spba=210.358n spba1=213.47n dfm_flag=0 sapb=217.823n
XM4 net305 eniob VDD VDD pch_12_mac l=70n w=12.0u multi=1 nf=12 sd=160.0n ad=9.6e-13 as=1.08e-12 pd=13.92u ps=16.16u nrd=0.003643 nrs=0.003643 sa=739.143n sb=739.143n sa1=320.464n sa2=597.542n sa3=827.446n sa4=691.15n sb1=320.464n sb2=597.542n sb3=827.446n spa=163.103n spa1=162.995n spa2=162.263n spa3=162.581n sap=276.12n spba=197.934n spba1=200.917n dfm_flag=0 sapb=299.055n
XM14 op headin net074 VDD pch_12_mac l=150.0n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM5 headin headin net071 VDD pch_12_mac l=150.0n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM13 on headref net068 VDD pch_12_mac l=150.0n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM12 headref headref net065 VDD pch_12_mac l=150.0n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM2 tailp vbiasp net305 VDD pch_12_mac l=200n w=16.0u multi=1 nf=16 sd=160.0n ad=1.28e-12 as=1.4e-12 pd=18.56u ps=20.8u nrd=0.002769 nrs=0.002769 sa=1.30442u sb=1.30442u sa1=377.952n sa2=893.294n sa3=1.06016u sa4=1.06817u sb1=377.952n sb2=893.294n sb3=1.06016u spa=160.613n spa1=160.608n spa2=160.565n spa3=160.593n sap=308.397n spba=248.146n spba1=255.744n dfm_flag=0 sapb=373.804n
XM24 on in net069 VDD pch_12_mac l=150.0n w=6u multi=1 nf=6 sd=160.0n ad=4.8e-13 as=6e-13 pd=6.96u ps=9.2u nrd=0.006918 nrs=0.006918 sa=532.241n sb=532.241n sa1=262.103n sa2=459.019n sa3=669.63n sa4=465.226n sb1=262.103n sb2=459.019n sb3=669.63n spa=161.639n spa1=161.625n spa2=161.519n spa3=161.582n sap=234.599n spba=225.543n spba1=231.605n dfm_flag=0 sapb=290.644n
XM18 op inb net085 VDD pch_12_mac l=150.0n w=6u multi=1 nf=6 sd=160.0n ad=4.8e-13 as=6e-13 pd=6.96u ps=9.2u nrd=0.006918 nrs=0.006918 sa=532.241n sb=532.241n sa1=262.103n sa2=459.019n sa3=669.63n sa4=465.226n sb1=262.103n sb2=459.019n sb3=669.63n spa=161.639n spa1=161.625n spa2=161.519n spa3=161.582n sap=234.599n spba=225.543n spba1=231.605n dfm_flag=0 sapb=290.644n
XM10 net065 eniob VDD VDD pch_12_mac l=70n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.009877 nrs=0.009877 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=202.288n spba1=205.319n dfm_flag=0 sapb=244.426n
XM7 net071 eniob VDD VDD pch_12_mac l=70n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.009877 nrs=0.009877 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=202.288n spba1=205.319n dfm_flag=0 sapb=244.426n
XM6 net074 eniob VDD VDD pch_12_mac l=70n w=4u multi=1 nf=4 sd=160.0n ad=3.2e-13 as=4.4e-13 pd=4.64u ps=6.88u nrd=0.009877 nrs=0.009877 sa=331.492n sb=331.492n sa1=220.515n sa2=312.483n sa3=477.658n sa4=315.144n sb1=220.515n sb2=312.483n sb3=477.658n spa=169.427n spa1=169.152n spa2=167.186n spa3=168.066n sap=217.368n spba=202.288n spba1=205.319n dfm_flag=0 sapb=244.426n
Xoffpin net069 offn12b[3] offn12b[2] offn12b[1] offn12b[0] eniob tailp VDD ckRxOffsetP
Xoffpinb net085 offp12b[3] offp12b[2] offp12b[1] offp12b[0] eniob tailp VDD ckRxOffsetP
.ends cmos12iAmpCore
.subckt sc_nand2x2l a b y inh_vdd inh_vss
XNb net21 b inh_vss inh_vss nch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.023481 nrs=0.023481 sa=201.53800n sb=201.53800n sca=2.27315 scb=0.000356871 scc=5.23214e-07 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XNa y a net21 inh_vss nch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.023481 nrs=0.023481 sa=201.53800n sb=201.53800n sca=2.27315 scb=0.000356871 scc=5.23214e-07 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XPb y b inh_vdd inh_vdd pch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
XPa y a inh_vdd inh_vdd pch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
.ends sc_nand2x2l
.subckt DamNcap2x2_12 minus plus
XC1 plus minus nmoscap_12 lr=2u wr=2u multi=1
.ends DamNcap2x2_12
.subckt ckRxLSBias en enb vbiasn vbiasp inh_vdd inh_vss
XM1 net26 enb inh_vdd inh_vdd pch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
XM0 vbiasp en inh_vdd inh_vdd pch_lvt_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
XP0 vbiasp vbiasp inh_vdd inh_vdd pch_lvt_mac l=150.0n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=230.068n sb=230.068n sca=10.4031 scb=0.00915566 scc=0.000801174 sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=179.221n spa1=178.832n spa2=175.961n spa3=177.655n sap=197.247n spba=235.815n spba1=242.211n enx=1.34301u enx1=1.33728u eny=383.886n eny1=216.004n eny2=305.235n rex=4.32095u rey=940.027n dfm_flag=0 sapb=244.813n sa5=235.841n sa6=331.192n sodx=140.0n sodx1=256.383n sodx2=883.875n sody=711.54n
XC0 inh_vss vbiasn DamNcap2x2_12
XXR5_1__dmy0 net26 XR5_1__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_2__dmy0 XR5_1__dmy0 XR5_2__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_3__dmy0 XR5_2__dmy0 XR5_3__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_4__dmy0 XR5_3__dmy0 XR5_4__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_5__dmy0 XR5_4__dmy0 XR5_5__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_6__dmy0 XR5_5__dmy0 XR5_6__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_7__dmy0 XR5_6__dmy0 XR5_7__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_8__dmy0 XR5_7__dmy0 XR5_8__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_9__dmy0 XR5_8__dmy0 XR5_9__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_10__dmy0 XR5_9__dmy0 XR5_10__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_11__dmy0 XR5_10__dmy0 XR5_11__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_12__dmy0 XR5_11__dmy0 XR5_12__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_13__dmy0 XR5_12__dmy0 XR5_13__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_14__dmy0 XR5_13__dmy0 XR5_14__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_15__dmy0 XR5_14__dmy0 XR5_15__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_16__dmy0 XR5_15__dmy0 XR5_16__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_17__dmy0 XR5_16__dmy0 XR5_17__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_18__dmy0 XR5_17__dmy0 XR5_18__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_19__dmy0 XR5_18__dmy0 XR5_19__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR5_20__dmy0 XR5_19__dmy0 vbiasn inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_1__dmy0 vbiasp XR4_1__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_2__dmy0 XR4_1__dmy0 XR4_2__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_3__dmy0 XR4_2__dmy0 XR4_3__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_4__dmy0 XR4_3__dmy0 XR4_4__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_5__dmy0 XR4_4__dmy0 XR4_5__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_6__dmy0 XR4_5__dmy0 XR4_6__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_7__dmy0 XR4_6__dmy0 XR4_7__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_8__dmy0 XR4_7__dmy0 XR4_8__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_9__dmy0 XR4_8__dmy0 XR4_9__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_10__dmy0 XR4_9__dmy0 XR4_10__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_11__dmy0 XR4_10__dmy0 XR4_11__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_12__dmy0 XR4_11__dmy0 XR4_12__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_13__dmy0 XR4_12__dmy0 XR4_13__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_14__dmy0 XR4_13__dmy0 XR4_14__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_15__dmy0 XR4_14__dmy0 XR4_15__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_16__dmy0 XR4_15__dmy0 XR4_16__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_17__dmy0 XR4_16__dmy0 XR4_17__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_18__dmy0 XR4_17__dmy0 XR4_18__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_19__dmy0 XR4_18__dmy0 XR4_19__dmy0 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XXR4_20__dmy0 XR4_19__dmy0 net29 inh_vss rppolywo_m lr=1.8u wr=1.8u multi=1 m=1
XM3 vbiasn enb inh_vss inh_vss nch_lvt_mac l=40n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=201.53800n sb=201.53800n sca=2.81171 scb=0.000664299 scc=1.04238e-06 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XM2 vbiasn vbiasn inh_vss inh_vss nch_lvt_mac l=150.0n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=230.068n sb=230.068n sca=2.76296 scb=0.000664288 scc=1.04238e-06 sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=179.221n spa1=178.832n spa2=175.961n spa3=177.655n sap=197.247n spba=235.815n spba1=242.211n enx=2.14718u enx1=2.14386u eny=1.00253u eny1=799.107n eny2=967.619n rex=4.18109u rey=1.86012u dfm_flag=0 sapb=244.813n sa5=235.841n sa6=331.192n sodx=140.0n sodx1=256.383n sodx2=883.875n sody=901.742n
XN0 net29 en inh_vss inh_vss nch_lvt_mac l=40n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=201.53800n sb=201.53800n sca=2.81171 scb=0.000664299 scc=1.04238e-06 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XM9 inh_vdd vbiasp inh_vdd inh_vdd pch_12_mac l=1u w=4.8u multi=1 nf=4 sd=160.0n ad=3.84e-13 as=5.28e-13 pd=5.44u ps=8.08u nrd=0.009075 nrs=0.009075 sa=982.244n sb=982.244n sa1=280.201n sa2=716.688n sa3=702.09n sa4=467.401n sb1=280.201n sb2=716.688n sb3=702.09n spa=162.463n spa1=162.444n spa2=162.362n spa3=162.458n sap=237.671n spba=305.922n spba1=367.073n dfm_flag=0 sapb=279.391n
.ends ckRxLSBias
.subckt sc_invx2r a y inh_vdd inh_vss
XP0 y a inh_vdd inh_vdd pch_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
XN0 y a inh_vss inh_vss nch_mac l=40n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=201.53800n sb=201.53800n sca=2.81171 scb=0.000664299 scc=1.04238e-06 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
.ends sc_invx2r
.subckt sc_nor2x2l a b y inh_vdd inh_vss
XNb y b inh_vss inh_vss nch_lvt_mac l=40n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=201.53800n sb=201.53800n sca=2.81171 scb=0.000664299 scc=1.04238e-06 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XNa y a inh_vss inh_vss nch_lvt_mac l=40n w=660.0n multi=1 nf=2 sd=160.0n ad=5.28e-14 as=9.24e-14 pd=980.0n ps=1.88u nrd=0.046963 nrs=0.046963 sa=201.53800n sb=201.53800n sca=2.81171 scb=0.000664299 scc=1.04238e-06 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=2.09649u enx1=2.09524u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.10544u rey=1.83014u dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=901.74200n
XPa y a net7 inh_vdd pch_lvt_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.7800n sb=309.7800n sca=10.2911 scb=0.00915362 scc=0.000801174 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=1.47532u enx1=1.46621u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.50641u rey=921.12900n dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=711.5400n
XPb net7 b inh_vdd inh_vdd pch_lvt_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.7800n sb=309.7800n sca=10.2911 scb=0.00915362 scc=0.000801174 sa1=217.49500n sa2=295.52600n sa3=447.84900n sa4=301.56200n sb1=217.49500n sb2=295.52600n sb3=447.84900n spa=169.42700n spa1=169.15200n spa2=167.14600n spa3=167.93300n sap=213.44600n spba=191.30700n spba1=193.11400n enx=1.47532u enx1=1.46621u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.50641u rey=921.12900n dfm_flag=0 sapb=245.13100n sa5=337.83200n sa6=438.67900n sodx=140.0n sodx1=304.44100n sodx2=947.8700n sody=711.5400n
.ends sc_nor2x2l
.subckt od12iLevelShift inn inp out outb rxen inh_vdd inh_vss
XM26 xn xn net065 inh_vss nch_lvt_mac l=150.0n w=1.2u multi=1 nf=2 sd=160.0n ad=9.6e-14 as=1.68e-13 pd=1.52u ps=2.96u nrd=0.021347 nrs=0.021347 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM28 xp xp net062 inh_vss nch_lvt_mac l=150.0n w=1.2u multi=1 nf=2 sd=160.0n ad=9.6e-14 as=1.68e-13 pd=1.52u ps=2.96u nrd=0.021347 nrs=0.021347 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM7 net065 xn inh_vss inh_vss nch_lvt_mac l=150.0n w=1.2u multi=1 nf=2 sd=160.0n ad=9.6e-14 as=1.68e-13 pd=1.52u ps=2.96u nrd=0.021347 nrs=0.021347 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM6 net062 xp inh_vss inh_vss nch_lvt_mac l=150.0n w=1.2u multi=1 nf=2 sd=160.0n ad=9.6e-14 as=1.68e-13 pd=1.52u ps=2.96u nrd=0.021347 nrs=0.021347 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM23 xn xp inh_vss inh_vss nch_lvt_mac l=40n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XM22 xp xn inh_vss inh_vss nch_lvt_mac l=40n w=300n multi=1 nf=1 sd=160.0n ad=4.2e-14 as=4.2e-14 pd=880.0n ps=880.0n nrd=0.068156 nrs=0.068156 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XM10 mirn inn net70 inh_vss nch_lvt_mac l=150.0n w=1u multi=1 nf=1 sd=160.0n ad=1.4e-13 as=1.4e-13 pd=2.28u ps=2.28u nrd=0.018546 nrs=0.018546 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM9 mirp inp net70 inh_vss nch_lvt_mac l=150.0n w=1u multi=1 nf=1 sd=160.0n ad=1.4e-13 as=1.4e-13 pd=2.28u ps=2.28u nrd=0.018546 nrs=0.018546 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM8 net70 vbiasn net113 inh_vss nch_lvt_mac l=150.0n w=2u multi=1 nf=4 sd=160.0n ad=1.6e-13 as=2.2e-13 pd=2.64u ps=3.88u nrd=0.018100 nrs=0.018100 sa=388.666n sb=388.666n sa1=227.236n sa2=354.562n sa3=541.173n sa4=345.184n sb1=227.236n sb2=354.562n sb3=541.173n spa=162.463n spa1=162.444n spa2=162.298n spa3=162.385n sap=212.983n spba=222.403n spba1=228.634n dfm_flag=0 sapb=266.153n
XM42 net113 en inh_vss inh_vss nch_lvt_mac l=40n w=16.0u multi=1 nf=16 sd=160.0n ad=1.28e-12 as=1.4e-12 pd=18.56u ps=20.8u nrd=0.001865 nrs=0.001865 sa=831.895n sb=831.895n sa1=346.58n sa2=654.425n sa3=889.782n sa4=800.916n sb1=346.58n sb2=654.425n sb3=889.782n spa=162.323n spa1=162.241n spa2=161.675n spa3=161.889n sap=287.862n spba=182.48n spba1=184.294n dfm_flag=0 sapb=279.467n
XM37 net112 enb inh_vdd inh_vdd pch_lvt_mac l=40n w=16.0u multi=1 nf=16 sd=160.0n ad=1.28e-12 as=1.4e-12 pd=18.56u ps=20.8u nrd=0.002769 nrs=0.002769 sa=831.895n sb=831.895n sa1=346.58n sa2=654.425n sa3=889.782n sa4=800.916n sb1=346.58n sb2=654.425n sb3=889.782n spa=162.323n spa1=162.241n spa2=161.675n spa3=161.889n sap=287.862n spba=182.48n spba1=184.294n dfm_flag=0 sapb=279.467n
XM35 tail vbiasp net112 inh_vdd pch_lvt_mac l=150.0n w=12.0u multi=1 nf=12 sd=160.0n ad=9.6e-13 as=1.08e-12 pd=13.92u ps=16.16u nrd=0.003643 nrs=0.003643 sa=919.751n sb=919.751n sa1=333.986n sa2=697.086n sa3=908.018n sa4=792.988n sb1=333.986n sb2=697.086n sb3=908.018n spa=160.818n spa1=160.811n spa2=160.753n spa3=160.787n sap=279.227n spba=229.023n spba1=234.869n dfm_flag=0 sapb=338.372n
XM16 xn mirn inh_vdd inh_vdd pch_lvt_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM15 mirn mirn inh_vdd inh_vdd pch_lvt_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM19 xp mirp inh_vdd inh_vdd pch_lvt_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM17 mirp mirp inh_vdd inh_vdd pch_lvt_mac l=150.0n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=170.0n spa1=170.0n spa2=170.0n spa3=170.0n sap=160.462n spba=201.742n spba1=208.507n dfm_flag=0 sapb=197.628n
XM34 xn inp tail inh_vdd pch_lvt_mac l=150.0n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM33 xp inn tail inh_vdd pch_lvt_mac l=150.0n w=2u multi=1 nf=2 sd=160.0n ad=1.6e-13 as=2.8e-13 pd=2.32u ps=4.56u nrd=0.017261 nrs=0.017261 sa=230.068n sb=230.068n sa1=177.935n sa2=223.401n sa3=331.644n sa4=213.865n sb1=177.935n sb2=223.401n sb3=331.644n spa=164.95n spa1=164.925n spa2=164.723n spa3=164.844n sap=182.796n spba=214.512n spba1=221.072n dfm_flag=0 sapb=229.376n
XM41 mirn en inh_vdd inh_vdd pch_lvt_mac l=40n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XM39 mirp en inh_vdd inh_vdd pch_lvt_mac l=40n w=500n multi=1 nf=1 sd=160.0n ad=7e-14 as=7e-14 pd=1.28u ps=1.28u nrd=0.075032 nrs=0.075032 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XU4 net067 out inh_vdd inh_vss sc_invx2l
XU3 net068 outb inh_vdd inh_vss sc_invx2l
XU6 crossn net068 inh_vdd inh_vss sc_invx2l
XU11 crossp net067 inh_vdd inh_vss sc_invx2l
XM27 crossp crossn net108 inh_vss nch_hvt_mac l=40n w=330.0n multi=1 nf=1 sd=160.0n ad=4.62e-14 as=4.62e-14 pd=940.0n ps=940.0n nrd=0.074972 nrs=0.074972 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XM43 crossn crossp net105 inh_vss nch_hvt_mac l=40n w=330.0n multi=1 nf=1 sd=160.0n ad=4.62e-14 as=4.62e-14 pd=940.0n ps=940.0n nrd=0.074972 nrs=0.074972 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XM31 net108 en inh_vss inh_vss nch_hvt_mac l=40n w=1.32u multi=1 nf=4 sd=160.0n ad=1.056e-13 as=1.452e-13 pd=1.96u ps=2.86u nrd=0.026879 nrs=0.026879 sa=309.78n sb=309.78n sa1=217.495n sa2=295.526n sa3=447.849n sa4=301.562n sb1=217.495n sb2=295.526n sb3=447.849n spa=169.427n spa1=169.152n spa2=167.146n spa3=167.933n sap=213.446n spba=187.09n spba1=188.941n dfm_flag=0 sapb=217.266n
XM38 net105 en inh_vss inh_vss nch_hvt_mac l=40n w=1.32u multi=1 nf=4 sd=160.0n ad=1.056e-13 as=1.452e-13 pd=1.96u ps=2.86u nrd=0.026879 nrs=0.026879 sa=309.78n sb=309.78n sa1=217.495n sa2=295.526n sa3=447.849n sa4=301.562n sb1=217.495n sb2=295.526n sb3=447.849n spa=169.427n spa1=169.152n spa2=167.146n spa3=167.933n sap=213.446n spba=187.09n spba1=188.941n dfm_flag=0 sapb=217.266n
XM30 net109 enb inh_vdd inh_vdd pch_hvt_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.78n sb=309.78n sa1=217.495n sa2=295.526n sa3=447.849n sa4=301.562n sb1=217.495n sb2=295.526n sb3=447.849n spa=169.427n spa1=169.152n spa2=167.146n spa3=167.933n sap=213.446n spba=187.09n spba1=188.941n dfm_flag=0 sapb=217.266n
XM32 net106 enb inh_vdd inh_vdd pch_hvt_mac l=40n w=2.64u multi=1 nf=4 sd=160.0n ad=2.112e-13 as=2.904e-13 pd=3.28u ps=4.84u nrd=0.019965 nrs=0.019965 sa=309.78n sb=309.78n sa1=217.495n sa2=295.526n sa3=447.849n sa4=301.562n sb1=217.495n sb2=295.526n sb3=447.849n spa=169.427n spa1=169.152n spa2=167.146n spa3=167.933n sap=213.446n spba=187.09n spba1=188.941n dfm_flag=0 sapb=217.266n
XM29 crossp crossn net109 inh_vdd pch_hvt_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.055711 nrs=0.055711 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XM44 crossn crossp net106 inh_vdd pch_hvt_mac l=40n w=660.0n multi=1 nf=1 sd=160.0n ad=9.24e-14 as=9.24e-14 pd=1.6u ps=1.6u nrd=0.055711 nrs=0.055711 sa=140.0n sb=140.0n sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.708n spba=191.625n spba1=193.742n dfm_flag=0 sapb=170.157n
XU5 xn en crossp inh_vdd inh_vss sc_nand2x2l
XI83 en enb vbiasn vbiasp inh_vdd inh_vss ckRxLSBias
XU1 enb en inh_vdd inh_vss sc_invx2r
XU0 rxen enb inh_vdd inh_vss sc_invx2r
XU15 xp enb crossn inh_vdd inh_vss sc_nor2x2l
.ends od12iLevelShift
.subckt DamNcap12 minus plus
XC1 plus minus nmoscap_12 lr=2u wr=2u multi=1
.ends DamNcap12
.subckt od12iAmp VDD in inb offcalen offtrim[4] offtrim[3] offtrim[2] offtrim[1] offtrim[0] out pd_rxen rxen inh_vdd inh_vss
XM46 xgateinp offcalenb in inh_vss nch_12_mac l=70n w=8u multi=1 nf=8 sd=160.0n ad=6.4e-13 as=7.6e-13 pd=9.28u ps=11.52u nrd=0.003584 nrs=0.003584 sa=545.317n sb=545.317n sa1=279.161n sa2=472.77n sa3=691.591n sa4=511.925n sb1=279.161n sb2=472.77n sb3=691.591n spa=164.669n spa1=164.513n spa2=163.442n spa3=163.91n sap=251.492n spba=198.962n spba1=201.956n dfm_flag=0 sapb=276.979n
XM0 xgateinn offcalenb inb inh_vss nch_12_mac l=70n w=8u multi=1 nf=8 sd=160.0n ad=6.4e-13 as=7.6e-13 pd=9.28u ps=11.52u nrd=0.003584 nrs=0.003584 sa=545.317n sb=545.317n sa1=279.161n sa2=472.77n sa3=691.591n sa4=511.925n sb1=279.161n sb2=472.77n sb3=691.591n spa=164.669n spa1=164.513n spa2=163.442n spa3=163.91n sap=251.492n spba=198.962n spba1=201.956n dfm_flag=0 sapb=276.979n
XM1 xgateinn offcalenbb inb VDD pch_12_mac l=70n w=16.0u multi=1 nf=16 sd=160.0n ad=1.28e-12 as=1.4e-12 pd=18.56u ps=20.8u nrd=0.002769 nrs=0.002769 sa=921.475n sb=921.475n sa1=353.378n sa2=702.745n sa3=930.644n sa4=860.283n sb1=353.378n sb2=702.745n sb3=930.644n spa=162.323n spa1=162.241n spa2=161.686n spa3=161.926n sap=295.864n spba=197.434n spba1=200.411n dfm_flag=0 sapb=316.19n
XM48 xgateinp offcalenbb in VDD pch_12_mac l=70n w=16.0u multi=1 nf=16 sd=160.0n ad=1.28e-12 as=1.4e-12 pd=18.56u ps=20.8u nrd=0.002769 nrs=0.002769 sa=921.475n sb=921.475n sa1=353.378n sa2=702.745n sa3=930.644n sa4=860.283n sb1=353.378n sb2=702.745n sb3=930.644n spa=162.323n spa1=162.241n spa2=161.686n spa3=161.926n sap=295.864n spba=197.434n spba1=200.411n dfm_flag=0 sapb=316.19n
XI81 VDD xgateinp xgateinn offcalen offcalenb offcalenbb offtrim[4] offtrim[3] offtrim[2] offtrim[1] offtrim[0] on op pd_rxen rxen inh_vdd inh_vss cmos12iAmpCore
XI84 on op out outb rxen inh_vdd inh_vss od12iLevelShift
XI80_10_ xgateinn inb DamNcap12
XI80_9_ xgateinn inb DamNcap12
XI80_8_ xgateinn inb DamNcap12
XI80_7_ xgateinn inb DamNcap12
XI80_6_ xgateinn inb DamNcap12
XI80_5_ xgateinn inb DamNcap12
XI80_4_ xgateinn inb DamNcap12
XI80_3_ xgateinn inb DamNcap12
XI80_2_ xgateinn inb DamNcap12
XI80_1_ xgateinn inb DamNcap12
XI80_0_ xgateinn inb DamNcap12
XI95_10_ xgateinp in DamNcap12
XI95_9_ xgateinp in DamNcap12
XI95_8_ xgateinp in DamNcap12
XI95_7_ xgateinp in DamNcap12
XI95_6_ xgateinp in DamNcap12
XI95_5_ xgateinp in DamNcap12
XI95_4_ xgateinp in DamNcap12
XI95_3_ xgateinp in DamNcap12
XI95_2_ xgateinp in DamNcap12
XI95_1_ xgateinp in DamNcap12
XI95_0_ xgateinp in DamNcap12
.ends od12iAmp
.subckt cxfr_12 D GN GP S inh_vdd inh_vss
XM1 S GN D inh_vss nch_12_mac l=70n w=4u multi=1 nf=8 sd=160.0n ad=3.2e-13 as=3.8e-13 pd=5.28u ps=6.52u nrd=0.009756 nrs=0.009756 sa=545.31700n sb=545.31700n sa1=279.16100n sa2=472.7700n sa3=691.59100n sa4=511.92500n sb1=279.16100n sb2=472.7700n sb3=691.59100n spa=164.66900n spa1=164.51300n spa2=163.44200n spa3=163.9100n sap=251.49200n spba=198.96200n spba1=201.95600n dfm_flag=0 sapb=276.97900n
XM5 S GP D inh_vdd pch_12_mac l=70n w=8u multi=1 nf=8 sd=160.0n ad=6.4e-13 as=7.6e-13 pd=9.28u ps=11.520u nrd=0.005323 nrs=0.005323 sa=545.31700n sb=545.31700n sca=4.26466 scb=0.00123141 scc=4.96875e-06 sa1=279.16100n sa2=472.7700n sa3=691.59100n sa4=511.92500n sb1=279.16100n sb2=472.7700n sb3=691.59100n spa=164.66900n spa1=164.51300n spa2=163.44200n spa3=163.9100n sap=251.49200n spba=198.96200n spba1=201.95600n enx=1.56827u enx1=1.51721u eny=520.0n eny1=520.0n eny2=520.0n rex=2.51924u rey=1.53982u dfm_flag=0 sapb=276.97900n sa5=600.14900n sa6=668.36100n sodx=490.0n sodx1=628.1800n sodx2=1.37524u sody=260.0n
.ends cxfr_12
.subckt sc_tiehilox1r tiehi tielo inh_vdd inh_vss
XN0 tielo tielo inh_vss inh_vss nch_mac l=40n w=330.0n multi=1 nf=1 sd=160.0n ad=4.62e-14 as=4.62e-14 pd=940.0n ps=940.0n nrd=0.074972 nrs=0.074972 sa=140.0n sb=140.0n sca=2.86377 scb=0.000664318 scc=1.04238e-06 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=2u enx1=2u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.0111u rey=1.83014u dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=901.74200n
XM0 tielo tiehi inh_vss inh_vss nch_mac l=40n w=330.0n multi=1 nf=1 sd=160.0n ad=4.62e-14 as=4.62e-14 pd=940.0n ps=940.0n nrd=0.074972 nrs=0.074972 sa=140.0n sb=140.0n sca=2.86377 scb=0.000664318 scc=1.04238e-06 sa1=140.0n sa2=140.0n sa3=140.0n sa4=140.0n sb1=140.0n sb2=140.0n sb3=140.0n spa=200n spa1=200n spa2=200n spa3=200n sap=178.70800n spba=221.26900n spba1=223.10500n enx=2u enx1=2u eny=977.48100n eny1=797.90800n eny2=967.61900n rex=4.0111u rey=1.83014u dfm_flag=0 sapb=210.88900n sa5=140.0n sa6=140.0n sodx=140.0n sodx1=206.67400n sodx2=831.18300n sody=901.74200n
XP0 tiehi tielo inh_vdd inh_vdd pch_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
.ends sc_tiehilox1r
XC0_5_ vref pwrn nmoscap_18 lr=2u wr=2u multi=1
XC0_4_ vref pwrn nmoscap_18 lr=2u wr=2u multi=1
XC0_3_ vref pwrn nmoscap_18 lr=2u wr=2u multi=1
XC0_2_ vref pwrn nmoscap_18 lr=2u wr=2u multi=1
XC0_1_ vref pwrn nmoscap_18 lr=2u wr=2u multi=1
XC0_0_ vref pwrn nmoscap_18 lr=2u wr=2u multi=1
XP0 offout rxenbb VREG VREG pch_mac l=40n w=1.32u multi=1 nf=2 sd=160.0n ad=1.056e-13 as=1.848e-13 pd=1.64u ps=3.2u nrd=0.034889 nrs=0.034889 sa=201.53800n sb=201.53800n sca=10.5905 scb=0.00916442 scc=0.000801174 sa1=173.19800n sa2=199.0600n sa3=267.47200n sa4=198.52500n sb1=173.19800n sb2=199.0600n sb3=267.47200n spa=179.22100n spa1=178.83200n spa2=175.72700n spa3=177.01700n sap=190.75200n spba=207.68900n spba1=209.41200n enx=1.2944u enx1=1.29231u eny=328.42100n eny1=214.58900n eny2=305.23500n rex=4.23096u rey=921.12900n dfm_flag=0 sapb=229.99700n sa5=211.51900n sa6=266.42600n sodx=140.0n sodx1=244.25600n sodx2=857.56100n sody=711.5400n
XI12 esel_odvref selbiasH selbiasL VDD VREG pwrn cmos12oLS
XI22 rxen net018 pd VDD VREG pwrn cmos12oLS
XU2 offout buf1 VREG pwrn sc_invx4r
XU5 buf2 rxoutB VREG pwrn sc_invx96r
XU4 buf1 buf2 VREG pwrn sc_invx20r
XU0 offout rxenbb rxenb lsout VREG pwrn cxfr m=1 nl=40n nw=330.0n nf=4 pl=40n pw=660.0n pf=4
XI5 vrefsel[0] vrefsel[1] vrefsel[2] vrefsel[3] vref pd VDD VREG pwrn vrefgen_error_in
XI9 pad VDD pwrn eEsdhbm
XI8 pad VDD pwrn eEsdhbm
XI11 pad in_esd VDD pwrn eEsdcdm
XI19 VDD in_esd vref net012 net012 net012 net012 net012 net012 lsout rxen rxen VREG pwrn od12iAmp
Xswibias emeas_odvref selbiasH selbiasL vref VDD pwrn cxfr_12
XI18_1_ net028[0] net012 VREG pwrn sc_tiehilox1r
XI18_0_ net028[1] net012 VREG pwrn sc_tiehilox1r
XU1 rxen rxenb VREG pwrn sc_invx1r
XU3 rxenb rxenbb VREG pwrn sc_invx1r
.ends od12i
